
library ieee;
use     ieee.std_logic_1164.all;


package pkg_OutputSamplesFi is

  type T_OUTPUTSAMPLESFI is array (0 to 2492-1) of std_logic_vector(35-1 downto 0);

  constant PKG_OUTPUTSAMPLESFI : T_OUTPUTSAMPLESFI := (
    "11111111110111101001100100111110010",
    "11111111110010001100111000111011001",
    "11111111110100111110011101011000110",
    "00000000000000101001010000011001011",
    "00000000001011111110100111000111111",
    "00000000001111100000100111000100110",
    "00000000001110011101010001011011010",
    "00000000001101110100010111100010000",
    "00000000001110101111100111101101110",
    "00000000001100010000100001101110101",
    "00000000000101100000101001000011010",
    "00000000000001000001110110101011111",
    "00000000000000101111010000010000111",
    "00000000000011001010111100001111101",
    "00000000000100100010001001101100110",
    "00000000000000100000001111001100100",
    "11111111111011000010001101110010010",
    "11111111111010111001101110010111010",
    "00000000000010010000100010001110110",
    "00000000001011110000101010110111111",
    "00000000010000111110000001000100100",
    "00000000010000001110100111111001100",
    "00000000001010111100101101101011111",
    "00000000000101001100110110110111001",
    "00000000000000000101110110011001000",
    "11111111111011110010011100110011001",
    "11111111111000101010001101010011000",
    "11111111110011010000011100111001111",
    "11111111101101110001011101010011101",
    "11111111101101111111010001111110011",
    "11111111110101100010001101010001011",
    "00000000000001011110100010110001010",
    "00000000001010001100010101100011001",
    "00000000001100001000111100111011010",
    "00000000000111100010100001001110010",
    "00000000000001110000000011001110000",
    "11111111111111000010000010100000011",
    "11111111111101010010011011011101100",
    "11111111111011110100110111110111000",
    "11111111111000001111110110010101001",
    "11111111110100100000111011011100011",
    "11111111110101110001000010010010010",
    "11111111111100101001010000111011001",
    "00000000000110011110011001000101001",
    "00000000001100111111101101111111000",
    "00000000001101100011000000101111100",
    "00000000001000111111010110111111001",
    "00000000000000111111100111100111010",
    "11111111111011101101101100100001000",
    "11111111111010111110001110101101100",
    "11111111111100011000110110100010010",
    "11111111111100011011101100100001111",
    "11111111111010010011011011011100001",
    "11111111111001011011000010100000101",
    "11111111111011001111001010011001100",
    "11111111111110000101010000010000000",
    "00000000000000110011100110000101110",
    "00000000000101001010110101010011100",
    "00000000001101010100011011011011011",
    "00000000010010110001111001001011010",
    "00000000001111010001010010100010000",
    "00000000000010101001101000010101010",
    "11111111110101110000010001100110101",
    "11111111110001101001101110111110001",
    "11111111110110000110111110010010001",
    "11111111111011111001001000000100100",
    "11111111111110111000101000010101011",
    "00000000000000100111111001001110100",
    "00000000000011101101011111101111110",
    "00000000000100111110101111100101111",
    "00000000000010010011000111000111000",
    "11111111111111010000110011000001000",
    "11111111111110110111101000110001100",
    "00000000000000100110100010010000000",
    "00000000000001100111001010010110100",
    "11111111111111101101111011101010011",
    "11111111111101111101001100110001000",
    "11111111111101001011010010100001110",
    "11111111111101000100001010111001101",
    "11111111111101110101011100101001111",
    "00000000000000111110011010001010100",
    "00000000000110000101100001100100101",
    "00000000001010000000011010110100110",
    "00000000001010010100101100000111001",
    "00000000000101000001011010001110000",
    "11111111111101011011110110000011100",
    "11111111111011001110100110111001001",
    "11111111111110101011010000001110100",
    "00000000000011001100101110111101010",
    "00000000000011010010010101110100010",
    "11111111111110000100011010111011100",
    "11111111111000110111000001000101010",
    "11111111110101111001101000000100000",
    "11111111110110111101000001100110110",
    "11111111111011000011101001101110001",
    "00000000000000111011010111110101100",
    "00000000000110001110101111100011111",
    "00000000000110101010101111111011111",
    "00000000000011100001011111110111011",
    "11111111111110100011010001001011011",
    "11111111111001110000010001010010100",
    "11111111111000100000101010111010100",
    "11111111111011110100100011001010111",
    "00000000000001010001110010111101000",
    "00000000000001000000101011101010001",
    "11111111111100001000110110101111001",
    "11111111111010000111111000110010010",
    "11111111111110101100001100001100010",
    "00000000000110010101010001011010101",
    "00000000001011011001001000111011001",
    "00000000001011011000111111101101101",
    "00000000000111101001101111001110101",
    "11111111111110101000010000110100000",
    "11111111110100000010011101001111110",
    "11111111110000010010001110110000101",
    "11111111110111111110101100000010001",
    "00000000000100001101100101101011001",
    "00000000001001110010011001001010111",
    "00000000000110100010111011100101001",
    "00000000000001110001000100001101001",
    "00000000000001111111101010000101111",
    "00000000000111111000100110110110101",
    "00000000001011011100010001111101111",
    "00000000001000001100111110010110110",
    "11111111111111001101100111110100101",
    "11111111110101101010111100100101001",
    "11111111101111101000100100101101110",
    "11111111101110011110000111111001010",
    "11111111110011010100101100100110100",
    "11111111111010000110111101100010101",
    "11111111111110110110000000111100110",
    "00000000000010011010111101001011010",
    "00000000000101011000000110110101001",
    "00000000001001011000000110100000100",
    "00000000001011101100001010110101010",
    "00000000001000100010111110011100010",
    "00000000000001001001100010111111011",
    "11111111111001000100001001000011000",
    "11111111110011111001110101110011111",
    "11111111110001000101011010000010010",
    "11111111110001001100101010101001001",
    "11111111110010011100001010110101000",
    "11111111110011001010010100100101010",
    "11111111110111010010100010111110101",
    "11111111111111011111111110100101110",
    "00000000001000010100101010001000000",
    "00000000001100100110011101100111110",
    "00000000001001100100011010111001011",
    "00000000000100000010000000010010010",
    "11111111111111010010000010110100010",
    "11111111111100000110000001111011100",
    "11111111111010001010001001101010101",
    "11111111111001010101110010101010111",
    "11111111111010001110111000110001110",
    "11111111111011110000000101100100010",
    "11111111111011010110001110101001000",
    "11111111111010101110000000101010101",
    "11111111111111001111111001110000110",
    "00000000001010001110100010100110010",
    "00000000010011101000110001111010011",
    "00000000010010110011011110000000011",
    "00000000000110100000111111111100111",
    "11111111111000011101111110011101011",
    "11111111110100010111000111011001100",
    "11111111110110111111010100001001010",
    "11111111110110000000111101110100111",
    "11111111110000100111110111111010100",
    "11111111101110000101001010011111010",
    "11111111110101100100010100111001001",
    "00000000000010101000111110011100110",
    "00000000001011111111001011001110000",
    "00000000001101000000101010101101110",
    "00000000001001000010010001001000110",
    "00000000000100101111010101100000000",
    "00000000000000010111000011011101101",
    "11111111111011100100001101110010101",
    "11111111110110111010011001110011100",
    "11111111110011001011111010011001011",
    "11111111110100100001001001000100011",
    "11111111111010000011101010011010010",
    "00000000000000000111111010101100110",
    "00000000000101011000011010011011000",
    "00000000001001011000011101001001110",
    "00000000001100000111001111111110010",
    "00000000001100010000000100010000100",
    "00000000001000000100001110000110001",
    "00000000000001010001100011111111010",
    "11111111111010111100110100111000010",
    "11111111110111100001100101011000111",
    "11111111110110110100101111100111000",
    "11111111111010010100011100011100000",
    "00000000000000010000001010011110101",
    "00000000000100001110100000101000010",
    "00000000000110011111101101000000010",
    "00000000000111001110010010111111100",
    "00000000000111001101111110100110000",
    "00000000000111100010111110011101101",
    "00000000000110110101100010010110101",
    "00000000000101100100100011110100001",
    "00000000000011111000100110000001001",
    "00000000000000100101001011000011101",
    "11111111111011100100110010110111100",
    "11111111110110111010101110110101100",
    "11111111110100100111010010010010111",
    "11111111110110001001011111101010001",
    "11111111111100110110011111110110110",
    "00000000000101001111010001011100110",
    "00000000001001100111000010101001011",
    "00000000001000100111100001110111100",
    "00000000000011101101100100101001100",
    "11111111111101110011000000001000010",
    "11111111111011000101011101011010000",
    "11111111111011110100010011111111100",
    "11111111111100101110010111010111100",
    "11111111111010110011110000001011011",
    "11111111111000010110111101111011100",
    "11111111111011011000000001100100110",
    "00000000000010001100101010111001000",
    "00000000000110100111011110000001000",
    "00000000000100100011010101110010110",
    "00000000000000101010000110101001001",
    "00000000000001101000110101100111101",
    "00000000000100101101100101000110011",
    "00000000000101111001011101001101110",
    "00000000000011101100010100110001101",
    "11111111111110110000011000001011001",
    "11111111111000011010111010011001001",
    "11111111110010000011000000101111000",
    "11111111101111110110011101000110011",
    "11111111110100011101110110001111000",
    "11111111111100000101101001010000101",
    "11111111111111010010001000101111000",
    "11111111111110000011000110100110011",
    "11111111111110010010001101101010000",
    "00000000000001100010100000111110100",
    "00000000000101011111110010010110100",
    "00000000000110001100101111111100011",
    "00000000000010100100101101100111010",
    "11111111111101111011011100010000100",
    "11111111111000010110011110000111100",
    "11111111110011000101101000011000010",
    "11111111110100001010111000110000111",
    "11111111111100010111010100110110001",
    "00000000000101101001000110000011010",
    "00000000001001011000101011110110100",
    "00000000000111010010110100001110100",
    "00000000000101010111101101110010000",
    "00000000000101111011111111001000000",
    "00000000000101000000011010000000010",
    "00000000000001101110101100100101000",
    "11111111111101011001010000110110011",
    "11111111111001110001000110010100001",
    "11111111111000001001100111001111100",
    "11111111111010111110011101110101001",
    "00000000000000101010100100110110110",
    "00000000000100101000110001010100001",
    "00000000000100010010011100000101001",
    "00000000000001101000110111011010101",
    "00000000000001111110000011011011100",
    "00000000000100101100101110001000001",
    "00000000000100000100011110101100011",
    "11111111111111001101101101000110010",
    "11111111111000111110000010001010100",
    "11111111110110010110101011000111110",
    "11111111110111000010001111101001010",
    "11111111111010100111011011001111101",
    "11111111111111111011011001011110101",
    "00000000000011111111000000111000001",
    "00000000000110001000000110011110011",
    "00000000000101100001000111100000010",
    "00000000000010110111110101101001010",
    "00000000000001111100101100100111111",
    "00000000000010100111010010011111101",
    "00000000000011010101011000111100010",
    "00000000000010011100001101000000000",
    "11111111111111100100111110111111111",
    "11111111111100100111101001110001100",
    "11111111111100000100100111011000011",
    "11111111111110111100101100000111100",
    "00000000000010100110011010010001101",
    "00000000000100000100110111111101011",
    "00000000000100000000011010001101100",
    "00000000000100000010001101000100000",
    "00000000000110011001000111001100111",
    "00000000000110101100000101001011010",
    "00000000000001011101010010101011100",
    "11111111111011010010100110101101100",
    "11111111111001010000101101101010001",
    "11111111111100111100101001001001111",
    "11111111111110011000111100110101010",
    "11111111111010010101101010000111110",
    "11111111110110001001101110111011101",
    "11111111110100001101101101101010001",
    "11111111110101101111111101110010011",
    "11111111111000000000100001111000000",
    "11111111111011000111111001010100000",
    "11111111111111111100000101001001110",
    "00000000000101011001100111010010101",
    "00000000001000100000000100001011100",
    "00000000000101110010001001100111100",
    "11111111111111101110110101101010110",
    "11111111111001110101011100110111001",
    "11111111110111000010110100101111111",
    "11111111111010000111001111011001111",
    "11111111111111110110110011111111001",
    "00000000000100000010010010111110010",
    "00000000000111010000110010101110111",
    "00000000001001011000111000101100111",
    "00000000001001100010101011010000100",
    "00000000000110000011011111100010001",
    "11111111111111000001110100110010001",
    "11111111111000011010100010001010010",
    "11111111110110010111000000110110001",
    "11111111111001100011110010100100011",
    "11111111111011100100110011010000100",
    "11111111111001111000000111111011111",
    "11111111110111110011001111010000110",
    "11111111111000001010111101111010001",
    "11111111111110001001111110010001001",
    "00000000000101100110000001111111101",
    "00000000001010000111000010100110000",
    "00000000001001001101101101000010001",
    "00000000000011100010000000011001101",
    "11111111111110001100100110110010101",
    "11111111111011010010011011011110011",
    "11111111111001110011011110011011110",
    "11111111110110111101010000111111100",
    "11111111110010100011111011111100100",
    "11111111101111111100110101001100000",
    "11111111110010000100110000000101111",
    "11111111111011110010000010000000101",
    "00000000001000000001001000010111110",
    "00000000001111000010100101010100001",
    "00000000001101000001111100100111011",
    "00000000000100100100011110010110110",
    "11111111111101000101000001010001011",
    "11111111111011001100011001100111011",
    "11111111111011100001111100011000001",
    "11111111111011011111100100011010011",
    "11111111111011110101111000000111101",
    "11111111111100010000101000111000000",
    "11111111111100110101000110101000101",
    "11111111111110100001101011001000011",
    "00000000000010001100110110100000101",
    "00000000000111011101010101011001100",
    "00000000001100110001111000001110101",
    "00000000001100111110011010000110001",
    "00000000000110011101001010001000011",
    "11111111111111110001011011100001001",
    "11111111111011111111111011000110001",
    "11111111111011010101010001111100100",
    "11111111111011111001010010110111001",
    "11111111111010111000111110010111110",
    "11111111111001101011000010101110110",
    "11111111111000110111111111101110011",
    "11111111111010001111100000111000011",
    "11111111111111010010001111000100111",
    "00000000000110010111100010010100001",
    "00000000001011100110011110110000011",
    "00000000001100011000110110100000010",
    "00000000001001001111011110110101000",
    "00000000000011100000101010111101001",
    "11111111111100100000000100101000000",
    "11111111110110011110110111100000111",
    "11111111110011000001111111000001110",
    "11111111110010110101110110000000011",
    "11111111110100011011101001011101011",
    "11111111110111111111110000100100010",
    "11111111111110001111110000100001100",
    "00000000000011101101000010100011110",
    "00000000000110101011001011110101011",
    "00000000000110111101101111011001110",
    "00000000000011000001001111001000011",
    "11111111111110100111110011011110010",
    "11111111111110110011101111001101011",
    "00000000000010100001101000100100110",
    "00000000000101010011001000000001011",
    "00000000000001011010001001010011011",
    "11111111111001101110001001011011101",
    "11111111110111010110101110101111000",
    "11111111111111000000111111000100011",
    "00000000001001110010010001110011101",
    "00000000001110110111011000001000001",
    "00000000001101010101100111100000111",
    "00000000001000000011100010100100110",
    "00000000000011011010010111001000001",
    "00000000000000001110110100001011100",
    "11111111111010111010011001001100101",
    "11111111110101100100110010001111001",
    "11111111110001100100001110100110010",
    "11111111110000000110111110100011100",
    "11111111110010000001111100011110011",
    "11111111110111001011111100101011001",
    "11111111111111000100101000110100100",
    "00000000000111100100010011110000001",
    "00000000001101010011100100010000110",
    "00000000001100111010011000000100001",
    "00000000000110000001011010000000100",
    "11111111111101001111011101100110100",
    "11111111110111100111110011110111001",
    "11111111110111011111000010001011011",
    "11111111111010001100100110000001101",
    "11111111111011101100100110111001111",
    "11111111111101001011011111000100000",
    "00000000000000111001101101000110101",
    "00000000000110001001011001001101101",
    "00000000001001000111011100111011001",
    "00000000000110010000011101001100000",
    "00000000000010010010101111010111000",
    "00000000000010000100011001010111100",
    "00000000000100011100111101000000101",
    "00000000000101001010010100011000000",
    "11111111111111111110101011000100010",
    "11111111110111111111111110101000101",
    "11111111110010000010011011101011000",
    "11111111110001000100100011010000010",
    "11111111110100011001011100110010100",
    "11111111111001111001111100110111101",
    "00000000000000001000101010100001001",
    "00000000000101100010111011100010000",
    "00000000001010000000101011010110010",
    "00000000001110011101101011010110001",
    "00000000010000001111010100011101001",
    "00000000001101101111001100110101000",
    "00000000000110100011111110110010101",
    "11111111111101101111111011001010010",
    "11111111111001011011011111110001101",
    "11111111111001110111000011000011001",
    "11111111111011000110100010011011010",
    "11111111111000100001010010001100000",
    "11111111110011100101111100101010111",
    "11111111110100110101000101000111001",
    "11111111111101110011110101001010100",
    "00000000001001010001010010100110000",
    "00000000001111001001111010000000100",
    "00000000001101001000011001000000101",
    "00000000000110110010100000111011100",
    "11111111111110010101010011110011011",
    "11111111110111111011111110001001101",
    "11111111110101000000011111100101110",
    "11111111110111011010100100101111110",
    "11111111111101111001110000100110000",
    "00000000000011001001001100101110100",
    "00000000000111011001010111000011111",
    "00000000001001101100000101000001111",
    "00000000000111110000001101100000010",
    "00000000000010111000101011110100101",
    "11111111111110101011011111100010010",
    "11111111111110100010100010010001100",
    "11111111111110011110101010010110011",
    "11111111111011011111011111110100110",
    "11111111110101110001000010011011001",
    "11111111110010010000110001100001110",
    "11111111110100001011011011001000000",
    "11111111111001100011001110100101111",
    "00000000000000001011000001010110100",
    "00000000000110111110100110010111110",
    "00000000001010100001101111001110111",
    "00000000001000111111110101100001100",
    "00000000000011011001000001011110000",
    "11111111111101010011101000001011001",
    "11111111111010100100100000001011110",
    "11111111111011011111101110100111111",
    "11111111111101010000101011101000111",
    "11111111111100101110000000101010010",
    "11111111111010100101111010001001010",
    "11111111111011001111010011111101110",
    "11111111111111000001111001010001110",
    "00000000000101010011011000100110010",
    "00000000001001011101011000000101001",
    "00000000001010000111010110100011011",
    "00000000001001011001111011101101101",
    "00000000000110110010010010100011001",
    "00000000000010101110011000100101110",
    "11111111111110000000110111001011001",
    "11111111111001011110110001111100011",
    "11111111110110001110010101110011010",
    "11111111110101111011111011100010010",
    "11111111111001100100111100110110100",
    "11111111111110100111110111100101110",
    "00000000000011000111110001100011111",
    "00000000000101100011001001011011100",
    "00000000000110100111110110100111111",
    "00000000001000011010100100111000110",
    "00000000001000101110101100110111110",
    "00000000000110001111011100111001001",
    "00000000000010000011001001000001101",
    "11111111111110101010010101110010100",
    "11111111111110011011100101110010001",
    "11111111111111010011010011111101100",
    "11111111111100101110000100110000000",
    "11111111110111001011100110100001100",
    "11111111110100100001101000110011011",
    "11111111111001101101000110001011111",
    "00000000000100001000100100111010111",
    "00000000001100011111011010111000111",
    "00000000001110100011000101010111100",
    "00000000001011010111011000101001010",
    "00000000000110111110100101111010101",
    "00000000000001011001101111100001101",
    "11111111111100111000001111110010010",
    "11111111111101110110110000000011111",
    "00000000000000011101110110000001110",
    "11111111111111001010101011000110011",
    "11111111111000110100110110111100000",
    "11111111110011010001001101101010101",
    "11111111110101001100101101111000101",
    "11111111111100110111011110100100000",
    "00000000000100001100100110010111101",
    "00000000000110110101101111011111000",
    "00000000000110010000111011100101100",
    "00000000000100011110100110101100111",
    "00000000000011110000110100011011111",
    "00000000000101011010101011000100111",
    "00000000000011010010001001111011001",
    "11111111111011101100111110001010101",
    "11111111110011111011101101100101010",
    "11111111110001100001111000000100000",
    "11111111110110001110100111000011101",
    "11111111111110011011010011101001001",
    "00000000000111001100100111110011110",
    "00000000001110001000110111011010100",
    "00000000001111001111001100101001110",
    "00000000001001010111111110000100100",
    "00000000000000110000010000001011101",
    "11111111111011111100010001100000001",
    "11111111111001110011100010101011100",
    "11111111110110111010111001101100111",
    "11111111110100110000110011110110011",
    "11111111110100101111101100010000100",
    "11111111110111011001110100100111110",
    "11111111111101001000001011000101101",
    "00000000000011010001101111110110100",
    "00000000001000011111001110000011100",
    "00000000001010001101100111110101001",
    "00000000001000001100010010100111001",
    "00000000000100100000000001100010110",
    "00000000000000100010000001100100111",
    "11111111111101011111010110111011111",
    "11111111111100000100011110111100001",
    "11111111111100110000000101010101010",
    "11111111111100110111101101101011011",
    "11111111111011000010001110001100101",
    "11111111111010101100010101011000111",
    "11111111111100111010110000100101010",
    "00000000000001100101011011110010010",
    "00000000000101110100011100110111011",
    "00000000000111101001100000011101001",
    "00000000000111001011011101010000001",
    "00000000000100010011100010001010010",
    "11111111111111110111000000100001100",
    "11111111111011001000010111111001101",
    "11111111111000001001111000010010100",
    "11111111111001001011100000001011100",
    "11111111111011110000110101010000010",
    "11111111111110100001000100001100001",
    "00000000000011010101101001000001011",
    "00000000001001101111001100110100010",
    "00000000001111001000010101110000110",
    "00000000001111010110010001101010101",
    "00000000001000111011100100001110001",
    "00000000000010101111100100000110001",
    "11111111111111111111110110010110111",
    "11111111111101100111101101101011001",
    "11111111111001111001110101011100111",
    "11111111111000001100100000010111100",
    "11111111111011101011101001101001001",
    "00000000000011001111000001011111010",
    "00000000001011010101101100001111110",
    "00000000001100110011101111101111101",
    "00000000000110101000100100111101101",
    "11111111111110111111000100001000010",
    "11111111111011000101101010111111011",
    "11111111111110100000011110010101011",
    "00000000000010111111101111110101111",
    "00000000000010001000011011100011100",
    "11111111111100111000100010111000110",
    "11111111110110100101100100000000001",
    "11111111110010101001001110001110010",
    "11111111110001111101011111101000101",
    "11111111110110101100011000111010111",
    "11111111111111010111000001011011001",
    "00000000000110001000100111110101010",
    "00000000001000001101101111111011111",
    "00000000000101001000011000100010101",
    "00000000000000101101101000111011000",
    "11111111111110000111110100010110100",
    "11111111111100100101001101000011100",
    "11111111111011111000001010101101001",
    "11111111111011101101100100000001001",
    "11111111111011110100101100011101101",
    "11111111111100110010000101010011101",
    "11111111111111100110100110001000010",
    "00000000000100011111001100010000010",
    "00000000001001111111001100111110000",
    "00000000001110111000101001110001010",
    "00000000001111111100111000110001111",
    "00000000001100101001101000001001110",
    "00000000001000100011011100100100100",
    "00000000000011111011100111111101000",
    "11111111111111000000100010011011101",
    "11111111111010101100111100010011100",
    "11111111111000000100100100110000101",
    "11111111111010001111010111110111100",
    "00000000000001000011111000111111101",
    "00000000000111001000000110110110110",
    "00000000001001110110001001001111010",
    "00000000001001000111111011111110001",
    "00000000000110001101010000011000010",
    "00000000000011011100110101011101111",
    "00000000000010010100011101101100010",
    "00000000000001100001101111010011110",
    "00000000000000010000111000100110111",
    "00000000000000100100101000101010001",
    "00000000000001100001101110011100110",
    "00000000000001110111011011100001111",
    "00000000000010101000011011111110100",
    "00000000000010101100100100011010011",
    "00000000000010010110010000111000110",
    "00000000000010001011010110101110000",
    "00000000000011001100000000000011001",
    "00000000000110110110110000000111010",
    "00000000001010001010111001011011111",
    "00000000001000011111100010010001000",
    "00000000000001101111100101011000110",
    "11111111111010110011100110011011110",
    "11111111110111010011000111000101000",
    "11111111110110000100000101110101111",
    "11111111110110100101011010111011101",
    "11111111111001000000110011111101000",
    "11111111111101001010100000101011011",
    "00000000000000100100000111001111011",
    "11111111111111011000001011111001010",
    "11111111111100011111011101000111110",
    "11111111111011000110100000010100001",
    "11111111111010001100100010000110011",
    "11111111111001001101111101001011010",
    "11111111110110001011011111111110000",
    "11111111110010010011101000010011011",
    "11111111110000111010011100100001010",
    "11111111110011011111110110111001010",
    "11111111111001010111011100000111000",
    "11111111111111110111001010011101011",
    "00000000000100010111001010111001100",
    "00000000000011111001001101010001111",
    "00000000000000110101101110010100100",
    "00000000000001111101001010010100100",
    "00000000000111101011100001111001111",
    "00000000001100001100000011011111110",
    "00000000000111101111000111011101010",
    "11111111111100001100111000110101001",
    "11111111110100001000101011110001111",
    "11111111110010110101010100001010011",
    "11111111110110111101111011001111111",
    "11111111111011111001011001101010000",
    "11111111111111001110011001010011000",
    "00000000000001011101000001011111111",
    "00000000000000101110101010111000001",
    "11111111111110110111011001010101010",
    "11111111111111011011001011101110010",
    "00000000000001111111001111001100110",
    "00000000000010001000110001111101000",
    "11111111111110001111110110011111110",
    "11111111111011101000010101110011000",
    "11111111111010110001101111110100100",
    "11111111111011001111001001010011011",
    "11111111111011101100011000001101011",
    "11111111111101011111010111000000111",
    "00000000000100100100000110110011100",
    "00000000001110100110111111100110010",
    "00000000010101111111011010001110000",
    "00000000010110010000111001010101111",
    "00000000001110100001010011010000101",
    "00000000000011110001000000000010111",
    "11111111111001111100010111000001010",
    "11111111110100011001010000000101011",
    "11111111110100000010110000010111001",
    "11111111110101111011100000101111001",
    "11111111110111011001000100001100001",
    "11111111110111110100100001011001011",
    "11111111111001111010100001011110000",
    "11111111111111000010100111011001110",
    "00000000000100100000101111010010111",
    "00000000000111001001100010100001000",
    "00000000000110110010001110011010101",
    "00000000000110100001101100000101101",
    "00000000000110110111011000010101010",
    "00000000000100010100110111100000001",
    "11111111111101000101101001111001101",
    "11111111110011110110111110111010011",
    "11111111101110110000100000011010100",
    "11111111110001101101001000111010100",
    "11111111111000110011101111010110001",
    "00000000000000000011001111001010100",
    "00000000000101100101011011111011110",
    "00000000001010001001100010010011011",
    "00000000001110011010111010010001000",
    "00000000001110001001010000011100001",
    "00000000001000100100101111110010110",
    "00000000000001110010100011001001001",
    "11111111111110001000110101011101110",
    "11111111111100011110001010100110101",
    "11111111111000010001010101011110100",
    "11111111110010100110101111001101100",
    "11111111101111001010110000011001110",
    "11111111110010011110110111010011011",
    "11111111111011100101010011111000011",
    "00000000000011000001101101101111001",
    "00000000000101011000101111001100000",
    "00000000000100010100110100100011110",
    "00000000000010110000000100001001111",
    "00000000000010111010001110011111011",
    "00000000000010000100110111100100100",
    "11111111111110010111100011101110010",
    "11111111111001010111011111000010101",
    "11111111110111100010111000001110111",
    "11111111111010001010111000110100111",
    "11111111111101111001010011001011000",
    "00000000000010000001101001101011011",
    "00000000000100111011100111111011001",
    "00000000000101000110101110101000110",
    "00000000000011111000100111011100010",
    "00000000000001110010000111011101111",
    "00000000000000111001101000011010011",
    "11111111111111100011001000000000001",
    "11111111111100100011011011110100110",
    "11111111110111011110011001010011011",
    "11111111110001000011110111000100000",
    "11111111101100110001111010110010101",
    "11111111101011110101111010100001100",
    "11111111101111011111100111101000101",
    "11111111110110111010100010100001111",
    "11111111111111000101110000001011101",
    "00000000000111001010111100110011010",
    "00000000001100110110111010010010100",
    "00000000001100110011100100111010011",
    "00000000000101011010101001101110011",
    "11111111111010000011111110001101111",
    "11111111110000111010011001111100000",
    "11111111101101111010100001000110110",
    "11111111110001110000111110100110001",
    "11111111111010001110011101100100100",
    "00000000000000011110010100110101011",
    "00000000000000101101001011000101110",
    "11111111111111101111011111011100000",
    "00000000000100111001010001111000100",
    "00000000001101111001010100111111100",
    "00000000010000101110111110110011000",
    "00000000001010111110011100001000101",
    "00000000000000111011111010011010001",
    "11111111111010011011110110110000010",
    "11111111111001100101000101101010011",
    "11111111110111111100011110100100111",
    "11111111110100011001000001110100101",
    "11111111110010101100001001001001101",
    "11111111110110001100001101000110001",
    "11111111111110100100100011101001111",
    "00000000000111011010100001011110111",
    "00000000001101001011100101101010111",
    "00000000001110010011100110111001000",
    "00000000001100001111111111001001011",
    "00000000000111111100010101110011001",
    "00000000000001111001011111011010010",
    "11111111111100001010001111110000010",
    "11111111110111000111000001000000011",
    "11111111110100000001110110111001000",
    "11111111110101011000010110001000001",
    "11111111111011000111000001110001100",
    "00000000000001000110101010111011100",
    "00000000000010010111110110010000001",
    "00000000000000100101011100000011110",
    "00000000000000101110000111110001111",
    "00000000000011011110000111001101110",
    "00000000000111100011011011111100111",
    "00000000001001010100110100100010000",
    "00000000000101110011011000011010000",
    "11111111111101100010011110110100110",
    "11111111110010100110101011110001011",
    "11111111101101101001100001001000000",
    "11111111110101000111100101000011011",
    "00000000000011101110110011100001111",
    "00000000001111000111101011000010011",
    "00000000010000110111011000010000000",
    "00000000001011010010000010101001100",
    "00000000000100001010011111100110110",
    "11111111111111100001000010010011011",
    "11111111111100010000001111111000000",
    "11111111111001101100000110101101001",
    "11111111111010000101010011101100000",
    "11111111111100110000110100010111011",
    "11111111111110111010001100001000100",
    "11111111111110011000100110011011110",
    "11111111111100001011101001110010001",
    "11111111111111101101010111000000101",
    "00000000001001001011110110000100001",
    "00000000001111101001001110100110001",
    "00000000001101000000000110110100011",
    "00000000000011110010001101000000111",
    "11111111111101011001100101100001010",
    "11111111111101010101100110110101001",
    "11111111111110101000111010101111011",
    "11111111111101011101000000000111110",
    "11111111111001001000110110111000010",
    "11111111110110011111000100110001101",
    "11111111110111101000001100101001001",
    "11111111111011010010100010110001110",
    "11111111111111011010010111110001101",
    "00000000000001111110101101110101101",
    "00000000000100001111100000010001101",
    "00000000000110101000101011110000100",
    "00000000000110111001111011000100000",
    "00000000000011001110001011101101000",
    "11111111111100111011001100100000011",
    "11111111111000100000100110100101001",
    "11111111110101110000001100111000000",
    "11111111110101100011100110100011011",
    "11111111110111010110110000010111001",
    "11111111111000100110111111001010101",
    "11111111111010111000011100010101111",
    "11111111111101011101100001111100110",
    "00000000000000010010111000011001111",
    "00000000000011011110100101100011110",
    "00000000000100010101100100010011110",
    "00000000000011010110110101111101000",
    "00000000000001100000110010100101010",
    "11111111111111010011011100001011110",
    "11111111111100110100111010100001000",
    "11111111111010100001101010100101011",
    "11111111111010110111010000011100101",
    "11111111111100110111111100101001100",
    "11111111111111110100010111011101111",
    "00000000000011100100001110111010101",
    "00000000000101010110011100100111110",
    "00000000000100111000111100101101101",
    "00000000000010110101001001110001100",
    "00000000000001111000101000000010000",
    "00000000000011000111000100011111000",
    "00000000000011100000011000100101100",
    "11111111111110011000101010000010110",
    "11111111110011011000101010000000110",
    "11111111101011101100000011100111010",
    "11111111101100111111101000100110010",
    "11111111110101110111011100011100010",
    "00000000000001001011101100011011000",
    "00000000000110000110110100001001111",
    "00000000000100010100110001111001010",
    "00000000000011101011000101100011011",
    "00000000000110110101001100111101111",
    "00000000001000001110111100101100010",
    "00000000000001101001111100110101000",
    "11111111110100101111100100101001111",
    "11111111101100011110100111000100000",
    "11111111101111111001101001100111111",
    "11111111111001100110111000100110101",
    "11111111111111110110100111010011110",
    "00000000000000111010011111110111110",
    "00000000000000110010000100110010101",
    "00000000000001011001001101000001101",
    "00000000000010001100001111000011110",
    "00000000000001010011000111111110111",
    "11111111111110110000111101001001011",
    "11111111111100001111011101000011110",
    "11111111111001001100001001111011001",
    "11111111110110011110011000011010110",
    "11111111110100001000100000001110000",
    "11111111110011000000000001001011010",
    "11111111110110001001000101000000000",
    "11111111111101110011101001011000111",
    "00000000000110111001000000000101001",
    "00000000001011001010101100111100011",
    "00000000000101111000101011110010111",
    "11111111111100100011110001110010101",
    "11111111111001010000101100100111001",
    "00000000000000000010000000010101100",
    "00000000001000010010001100010011111",
    "00000000000111001000100000101100010",
    "11111111111011101100100010000010111",
    "11111111110001101110001011001101110",
    "11111111110011100001101110110111010",
    "11111111111011101111010001110110111",
    "00000000000001011000110000011001000",
    "00000000000001111100011010101100000",
    "11111111111111111000100011011001010",
    "11111111111111110101011011011010011",
    "00000000000010010011010101110010010",
    "00000000000101001101100001110100010",
    "00000000000111010101111001110011000",
    "00000000000101110000111101000101111",
    "11111111111111010101011110010100100",
    "11111111110110110001011111010010110",
    "11111111110000010010010100000011001",
    "11111111110000100111000001011110101",
    "11111111110111110110011110011001001",
    "00000000000010000100000000111011110",
    "00000000001001010111001111110100110",
    "00000000001010000010110111010100000",
    "00000000000111110000100010011010011",
    "00000000000110110010111101010010000",
    "00000000000111110011010101111101111",
    "00000000000100111110101100011000010",
    "11111111111100111100100111111000010",
    "11111111110100111111001110000010100",
    "11111111110001000110010111001001000",
    "11111111110010100100100111011000010",
    "11111111110110111001000100100101100",
    "11111111111101000111110001101010110",
    "00000000000101101101010110011111010",
    "00000000001011101001110111011010100",
    "00000000001010101111001111111111001",
    "00000000000011001100011111101011100",
    "11111111111010100000100001001010010",
    "11111111110101100011110001101111001",
    "11111111110100010010000011111101110",
    "11111111110111111000001010001001110",
    "11111111111110011111101101100011011",
    "00000000000011000011111000100000001",
    "00000000000011000000010000111010000",
    "11111111111111111101010011111100000",
    "00000000000000011101101100000011010",
    "00000000000110100111101100110110010",
    "00000000001101001110100010111010101",
    "00000000001110000011111001100100100",
    "00000000001000111100110010111111000",
    "00000000000011010011000100110011111",
    "11111111111101101111100011001110011",
    "11111111111000111110101010011000010",
    "11111111110111001100000111010010101",
    "11111111110110110001011011000010111",
    "11111111110110011100001111010010010",
    "11111111110110111000110100010110001",
    "11111111111010111110110011000100101",
    "00000000000100101110110101010001000",
    "00000000001100111011110110110011000",
    "00000000001101110100000010101111001",
    "00000000001001010001100010000010001",
    "00000000000110101101010110010000000",
    "00000000000110010000100111011101110",
    "00000000000010001111010100011011100",
    "11111111111100011001010001101000010",
    "11111111111000100001110100010100001",
    "11111111110111111011100110110000110",
    "11111111111001000101100011101110101",
    "11111111111001111100111110011010110",
    "11111111111101001010000111101101011",
    "00000000000010101010111011001001110",
    "00000000000111010101100001000010011",
    "00000000000111001101011000100111000",
    "00000000000010100011101110101111011",
    "11111111111111101100111011101011011",
    "11111111111111011010111001000100110",
    "11111111111111010010011001111111101",
    "11111111111110111101011010100100001",
    "11111111111111011101001000101100011",
    "00000000000010010000101111010001000",
    "00000000000011111001111000010110110",
    "00000000000010100010001011001010000",
    "00000000000001011000111010101010100",
    "00000000000010101111010001110010000",
    "00000000000101111000010110001000100",
    "00000000000110011101010110000011111",
    "00000000000101100011000001000111001",
    "00000000000101100000010101110011110",
    "00000000000100101110011001100000110",
    "00000000000000101111011011100011110",
    "11111111111010011001110100101110010",
    "11111111110110000111101011001110100",
    "11111111110110011100111101111101111",
    "11111111111011001010101100100010110",
    "00000000000011001001101100110010101",
    "00000000001001111010101100010000100",
    "00000000001011011001100111111000110",
    "00000000001010011100110011110011111",
    "00000000001011101110100101110010110",
    "00000000001101110010010101011101010",
    "00000000001010011110001111001000001",
    "00000000000001101110001011100101110",
    "11111111111001011111111001100110111",
    "11111111110111000001101100100101100",
    "11111111111011110110110110110101110",
    "00000000000010110000100110110101001",
    "00000000000111111101110000000101100",
    "00000000001011010000111111110011000",
    "00000000001000110111101110000101011",
    "00000000000010100100001001000110001",
    "11111111111101010000111111100111101",
    "11111111111010110011110000001100110",
    "11111111111001111010100111100001101",
    "11111111111001010111100110111001001",
    "11111111111010101010101100001001000",
    "11111111111110001100010010001011011",
    "00000000000001010010110101001011001",
    "00000000000010100111001101011110101",
    "00000000000001101101111101001100111",
    "00000000000001111110110111101001111",
    "00000000000100011010010110011111010",
    "00000000000111010010100100000000000",
    "00000000000111001110010000000110101",
    "00000000000100010001010100100110011",
    "00000000000001110010011110000001100",
    "11111111111110011011001010111100000",
    "11111111111001110100011110110101000",
    "11111111110101110110011011101001011",
    "11111111110011110001100100001100110",
    "11111111110110000100110011000101111",
    "11111111111011110001000010100010000",
    "00000000000000011011010100000100101",
    "00000000000000100010010111110000011",
    "11111111111110110011101101010100011",
    "00000000000001001001001001100010000",
    "00000000001000100001111100100000010",
    "00000000001111011001111110111001100",
    "00000000001110011111000000011101100",
    "00000000000101001000011111110010000",
    "11111111111100000100100001111001010",
    "11111111111000011010011011000000011",
    "11111111110111100101101011111101001",
    "11111111111000000000000001111010110",
    "11111111111000101110110001100000010",
    "11111111111010110101001101111011101",
    "00000000000000110111100000011000000",
    "00000000001001110101101111000111100",
    "00000000010000111110100110001000000",
    "00000000001111010101011001100001001",
    "00000000000101010011101111000101001",
    "11111111111011110110001001101011100",
    "11111111111001000111100000101111101",
    "11111111111011101011001110111111100",
    "11111111111100101001011000000011010",
    "11111111111010111010001001101010001",
    "11111111111010011010111111110100100",
    "11111111111101000101101110011110001",
    "00000000000010011111011111001110010",
    "00000000001001010100110010000110110",
    "00000000010011011001101011100110001",
    "00000000011001101100111100101111010",
    "00000000010100011110101110100000111",
    "00000000000110101001010110000010101",
    "11111111110111101110111001000110010",
    "11111111110000001000111100101110011",
    "11111111101110011100000101001010110",
    "11111111101111110111010110101011111",
    "11111111110101111001000001110111101",
    "11111111111110011101100101000000010",
    "00000000000101000011011001011101101",
    "00000000000111011011101101011101111",
    "00000000001001000110001110101001011",
    "00000000001100100011010110001011101",
    "00000000001111001110011101010000111",
    "00000000001101011100101101001011000",
    "00000000000111001001101101111101001",
    "00000000000000101000010010101100111",
    "11111111111010110111011001111111011",
    "11111111110101111000110001011001100",
    "11111111110101000010010111011101110",
    "11111111111000011001001011000101011",
    "11111111111101011101000110010111010",
    "00000000000010111111100001011101010",
    "00000000000111101010100000110000000",
    "00000000001011010110111010010110000",
    "00000000001100111011101011000100100",
    "00000000001011001001011100101111000",
    "00000000000101101011110000010111011",
    "11111111111101110100110000001010100",
    "11111111111000101110101111100001100",
    "11111111110111100010001110000110110",
    "11111111111010000000010100110011111",
    "11111111111111010001001101010010111",
    "00000000000011111100111011100001101",
    "00000000000110110011111011010111000",
    "00000000000111000111010000110000010",
    "00000000000100101110100110010010011",
    "00000000000000101000000100001001000",
    "11111111111110010011011010111001101",
    "00000000000000001101100100010010101",
    "00000000000010110001011101000110010",
    "00000000000100111111001001111000000",
    "00000000000100011011010001101110011",
    "11111111111110100011100111010101111",
    "11111111110111000110100100100101011",
    "11111111110100101000110010111100000",
    "11111111111010000010011100111100011",
    "00000000000010010110100001100000001",
    "00000000000110001011010101010111000",
    "00000000000100110101111011000100011",
    "00000000000011111011100110011111101",
    "00000000000110011100010000011111100",
    "00000000000101110000111001100111001",
    "11111111111101010010010000001000101",
    "11111111110011011101000100110101011",
    "11111111110010010010000010010001000",
    "11111111111010011111010011000101000",
    "00000000000011001101111110011011010",
    "00000000000011000001110111100100010",
    "11111111111100011100111100010111010",
    "11111111111000010000111111110000001",
    "11111111111100001011010100111010000",
    "00000000000101010011000110110010010",
    "00000000001001010111101011001111110",
    "00000000000011111011011101010001011",
    "11111111111010100111010100000100101",
    "11111111110101111111110110010011110",
    "11111111110111100101001101001110011",
    "11111111111001011110111011011001101",
    "11111111110111110100111000001100110",
    "11111111110011111001001110001000001",
    "11111111110100110011001111001101000",
    "11111111111101010001110101000010000",
    "00000000000110110100111100110111100",
    "00000000001010111111001001000101111",
    "00000000000110101000100101110010010",
    "11111111111110010110011001001110010",
    "11111111111011100010010111000111000",
    "11111111111110110101010100011110001",
    "00000000000010101010111111100100110",
    "00000000000001111110111100000001011",
    "11111111111101000100101110001101010",
    "11111111111000101101111101011111101",
    "11111111111001001010110000111000010",
    "00000000000000110001011100100000100",
    "00000000001011010101100010101110110",
    "00000000010010000011000010010000011",
    "00000000010001001001110000011001001",
    "00000000001010001111111110111101110",
    "00000000000011100111011001010001000",
    "11111111111110011100000101100111100",
    "11111111111011010111001110011010010",
    "11111111111010111001110011011110000",
    "11111111111010111100001001011011000",
    "11111111111100010100000101001100001",
    "11111111111110100001101111111000111",
    "00000000000000010010011010111100111",
    "00000000000010110110010010011011110",
    "00000000000110011110110010101111011",
    "00000000001010111001110110011100100",
    "00000000001100111011100110111100011",
    "00000000001010010000000101000100110",
    "00000000000011111010100000011000110",
    "11111111111101110001010011111000111",
    "11111111111010100111010111011100011",
    "11111111111000000001111001010011000",
    "11111111110110111000001001111101110",
    "11111111111001110100100011010000100",
    "00000000000001000010010001101010111",
    "00000000001001101100000011001110101",
    "00000000001101000000000001000111111",
    "00000000001001101010100000000101101",
    "00000000000101001000100000010011101",
    "00000000000001100101001111110001011",
    "11111111111110101010010010110101011",
    "11111111111011010000100111101100000",
    "11111111111000100111001111010101100",
    "11111111111001100001011000011111001",
    "11111111111100011000010100010111011",
    "11111111111100110111000000000111111",
    "11111111111011000101001000110010001",
    "11111111111010110010110001100110011",
    "11111111111100110100000111101110100",
    "00000000000001000000111001110000011",
    "00000000000111111100110000100110111",
    "00000000001110000100010010111101111",
    "00000000001110001110010110110101000",
    "00000000001000001110101000100101111",
    "11111111111111011000010111111110101",
    "11111111111001101010011001110100000",
    "11111111110111100011010100100101100",
    "11111111110110011101111001010011000",
    "11111111110111010011101000101101110",
    "11111111111001110000000111101010101",
    "11111111111111011001100101001001001",
    "00000000000111110011000111110001010",
    "00000000001101101010100110110100000",
    "00000000001111111101100010000110000",
    "00000000001110000101111010010101000",
    "00000000001010101010110000111110110",
    "00000000000101001101000000001001011",
    "11111111111101111111100000110001000",
    "11111111110111011000100010011101010",
    "11111111110101001111011110110100010",
    "11111111111001111100100001111001001",
    "11111111111110011100011110000110100",
    "00000000000001110110101001100001100",
    "00000000000110111100011111011101000",
    "00000000001001010000010100000001100",
    "00000000000110111000010111110110010",
    "00000000000000111101011001111110110",
    "11111111111101010001100000100011111",
    "11111111111101011110101100101111001",
    "11111111111100001000110001001111000",
    "11111111110110100010001110001101001",
    "11111111110000101010011001000010110",
    "11111111101111111110010010100101001",
    "11111111110011100111000111000100010",
    "11111111110110111100110100011010100",
    "11111111111010111000011110101000101",
    "11111111111111100010001010001101000",
    "00000000000101001010111000100010110",
    "00000000001011000001111011010101100",
    "00000000001100111100000101100001100",
    "00000000001000001100000100000110110",
    "11111111111101111000101100011011111",
    "11111111110101100111010000001001100",
    "11111111110101001101110011010100111",
    "11111111111001111011000101011110100",
    "11111111111111011101100111001010111",
    "00000000000001011010000010000000001",
    "00000000000001111000001010100110111",
    "00000000000010000101100000001000100",
    "11111111111111110010001100101110100",
    "11111111111101001111110000001101000",
    "11111111111101010101110010001001000",
    "00000000000001101100110100100101001",
    "00000000001000110001001111111101010",
    "00000000001010100001001110110111110",
    "00000000000011011000100111000110100",
    "11111111111001010011101001101011011",
    "11111111110101111000010100010101111",
    "11111111111010010110110110100100011",
    "00000000000000100100000100000011000",
    "00000000000100010100010000101110110",
    "00000000000110010101001100010101001",
    "00000000001010001111100011111000001",
    "00000000001101100000011010111010111",
    "00000000001011010100110101001011101",
    "00000000000101011010110010011111100",
    "11111111111110111000010101011010010",
    "11111111111010010100000111101001001",
    "11111111111001110110110111110010101",
    "11111111111011110011000101110110101",
    "11111111111101000000110100111001010",
    "11111111111011100110101010111001010",
    "11111111111001011110011110100000101",
    "11111111111011010111100111010110110",
    "00000000000001110000111001110111011",
    "00000000001010011111111100101110010",
    "00000000001111111010110111000110001",
    "00000000001100101001101110110100101",
    "00000000000010111001101111110100111",
    "11111111110111110000110001010010111",
    "11111111110010000000001000011100111",
    "11111111110100001111000100010111010",
    "11111111111010101010101011011111001",
    "11111111111111111000000111010011111",
    "00000000000010001011001100010001110",
    "00000000000100101100111010011010101",
    "00000000001000011100110010111110100",
    "00000000001101100111001010100001001",
    "00000000010001100010101101011001101",
    "00000000010000011000110101111011111",
    "00000000001100010001110111000000010",
    "00000000000110010110001010110100101",
    "11111111111111001110111110000101101",
    "11111111111010000001110010001010010",
    "11111111110110101001011100111110110",
    "11111111110110011010111000000010110",
    "11111111111001100010110101101111111",
    "00000000000000011100000110100101010",
    "00000000001001110111100010110000000",
    "00000000010000011100101111101101110",
    "00000000010000110101101000100001011",
    "00000000001101101101111000010100111",
    "00000000001101011110101010101110011",
    "00000000001110101010010010111111000",
    "00000000001011001110111010010101000",
    "00000000000010010110100111000101110",
    "11111111110111101000101110000010100",
    "11111111110001110000011011110001001",
    "11111111110010101101111111000111000",
    "11111111111001011100101100001001010",
    "00000000000100000001101111000101000",
    "00000000001101110100100100011001100",
    "00000000010001010001100111011001001",
    "00000000001101110001100100010000000",
    "00000000001000101000000010010111111",
    "00000000000110111110000100011011001",
    "00000000000111001000011100110010101",
    "00000000000011111010110010011001001",
    "11111111111100100000001011011000101",
    "11111111110100111001100000001000111",
    "11111111110101010110111101101001101",
    "11111111111110111111111101111011001",
    "00000000001001111011001011011101010",
    "00000000001110000011111101011100000",
    "00000000001011001101110111101001010",
    "00000000001000101001010011000010010",
    "00000000001000000000011110100100011",
    "00000000000111001001000010010010101",
    "00000000000101001101110111100000011",
    "00000000000011011111100000100000010",
    "00000000000010111010011010011101010",
    "11111111111111111110111110010100110",
    "11111111111011001111000011111011000",
    "11111111111000111000101011000111100",
    "11111111111011001100011110000111100",
    "11111111111111010010110000000110010",
    "00000000000010000100010111110000101",
    "00000000000011111000010101100101100",
    "00000000000100111111001010011011011",
    "00000000000101101111010010000101111",
    "00000000000110101110110010110100001",
    "00000000000110011101111100001101000",
    "00000000000010110000100010101111010",
    "11111111111100110000000011110001000",
    "11111111111000101110110101011100010",
    "11111111111011001101111101001101001",
    "00000000000001001100111110000001000",
    "00000000000100000011000011011111010",
    "00000000000011010101000100011001110",
    "00000000000011010100011111111100000",
    "00000000001000010111000000111101100",
    "00000000001110001010101101101111000",
    "00000000001101111110110100001010001",
    "00000000000110111110000111001111111",
    "11111111111101011101101101001010010",
    "11111111111000001110101100100001000",
    "11111111110110111111111110001110001",
    "11111111110110100011011100010001001",
    "11111111110110010011101010000111011",
    "11111111110111011000110011111000001",
    "11111111111011000110110111110111100",
    "00000000000000000110000000000001010",
    "00000000000101010100100111111010111",
    "00000000001000110001100110001101010",
    "00000000000111111011101111011010010",
    "00000000000011110001001101111000001",
    "11111111111110111110100100001001000",
    "11111111111101010001101011000001100",
    "11111111111110001010101000011001111",
    "11111111111110001101000010001111101",
    "11111111111110001001010111000010101",
    "11111111111110111100011010001001101",
    "11111111111111100111010010001100100",
    "11111111111101110011101100110100100",
    "11111111111001011011100101111001011",
    "11111111110111111011110011101100101",
    "11111111111011001010011111000110100",
    "11111111111111011100011100110001100",
    "00000000000000010010011100001111001",
    "11111111111100000111110010001111001",
    "11111111110110110010111110001101100",
    "11111111110011001100010011100100011",
    "11111111110100100111110001100011001",
    "11111111111100101001000010110010100",
    "00000000000110110110000111010010010",
    "00000000001101000011101101010110001",
    "00000000001011111110110001101010010",
    "00000000001000010000001111110110111",
    "00000000000101111001111111011101111",
    "00000000000010111010010010110100010",
    "11111111111110110110011001001010100",
    "11111111111010100011111001100111010",
    "11111111111000001011111100001100110",
    "11111111111000000001101011010101011",
    "11111111111000111101110110001110001",
    "11111111111101001011111001011110111",
    "00000000000011001100111010000110111",
    "00000000000101010110101111110111011",
    "00000000000001111110010011100111010",
    "11111111111110111110011100111010011",
    "00000000000010011100010011011101100",
    "00000000001000000111011101110110011",
    "00000000001001111111000100110101010",
    "00000000000111100000010111110101111",
    "00000000000011000111111000110001110",
    "11111111111111000001100100000010110",
    "11111111111001001010010101100000101",
    "11111111110100001101000011011101000",
    "11111111110101010101100001001000101",
    "11111111111100000111101100001001100",
    "00000000000100110011110111110100100",
    "00000000001010001110000010110000011",
    "00000000001011000100101110100001001",
    "00000000001001111101101000001011100",
    "00000000000111010001101000100101100",
    "00000000000010110010101111111000111",
    "11111111111101000101000000001011011",
    "11111111111000011111111010010000001",
    "11111111110111100100010100110001010",
    "11111111111010011111010101111110101",
    "11111111111111010010001001100011101",
    "00000000000010000001110111001010100",
    "00000000000010010100111011111111011",
    "00000000000010001101100001101100100",
    "00000000000011001000110110110100100",
    "00000000000110110001010111010011001",
    "00000000001001000110010110011110000",
    "00000000000111100010110101000010011",
    "00000000000101001000101011010001110",
    "00000000000100001101001100001110010",
    "00000000000100011011011001111111010",
    "00000000000001011100010000100000010",
    "11111111111010111000100011010000000",
    "11111111110111001100111010000010000",
    "11111111111001101101110111011000100",
    "11111111111110000101100110000101100",
    "11111111111111101000110010101111110",
    "11111111111110110101101100001001101",
    "00000000000001011001000000110100110",
    "00000000000110101111011001011110010",
    "00000000001000011100010000010010111",
    "00000000000011000111111000110101111",
    "11111111111010110001010110011011110",
    "11111111110110000010011001011000000",
    "11111111110100110011011100001101100",
    "11111111110110001000110011101100010",
    "11111111111001111101011000110010110",
    "00000000000000001100001001101010011",
    "00000000000101010100111011111100111",
    "00000000000010100001010011000101010",
    "11111111111100110011000000111110000",
    "11111111111011101011101011100000001",
    "00000000000000100001111111111010110",
    "00000000000110010100111100110000110",
    "00000000000100100001001010111100010",
    "11111111111101011111101010110001000",
    "11111111110111111001111010111110110",
    "11111111110110110111100000011110010",
    "11111111111000110100111101110101000",
    "11111111111100001010000111001101011",
    "11111111111111100001101110101110101",
    "00000000000000111001110100111001110",
    "00000000000001110101011110001111010",
    "00000000000100110010111111101101111",
    "00000000001001101110111000111011010",
    "00000000001111011001110001100010100",
    "00000000001111100100110001100100110",
    "00000000000110110101100101010010010",
    "11111111111001011001000100011110100",
    "11111111101110100111001100100100011",
    "11111111101101111101001110010011000",
    "11111111110110100001011000010111100",
    "00000000000000010000111110111000000",
    "00000000000110110000100010011001001",
    "00000000001000100000011101101000010",
    "00000000001000010110001111101010101",
    "00000000000111110010000011010110110",
    "00000000000101101000101000000100110",
    "00000000000010100110010011111001010",
    "00000000000000011010011011100110011",
    "00000000000000001001010100111011001",
    "11111111111111000111100000111010001",
    "11111111111101001100011001110101011",
    "11111111111011101110011111000101010",
    "11111111111100100000010000100111010",
    "00000000000001101100000111001110011",
    "00000000000110100001101010000001110",
    "00000000000110011001101110001100110",
    "00000000000100111001111001000011100",
    "00000000000101111000011011001111000",
    "00000000001000011100001011001101101",
    "00000000000110101101101011011101010",
    "11111111111110100110011001100101010",
    "11111111110101001101010010010110001",
    "11111111110000111110110100011010100",
    "11111111110100011000101110011010010",
    "11111111111010100000111111101011001",
    "11111111111111101010011011001101100",
    "00000000000011001100111111010010001",
    "00000000000011110110000111111101011",
    "00000000000010100011000111000011100",
    "00000000000000001110000111001100110",
    "11111111111101011001001001011111010",
    "11111111111010010110001010000000001",
    "11111111110111010000010100001011110",
    "11111111110100101111100011011101110",
    "11111111110010010111101110010110011",
    "11111111110010001100100111011111100",
    "11111111110101000010000101011111001",
    "11111111111010010011100100111100111",
    "00000000000000111010010110010000111",
    "00000000000101110100100101101011001",
    "00000000000110100100011101010010100",
    "00000000000100010101110000010101000",
    "00000000000000011110011110110111111",
    "11111111111100100110100100101111101",
    "11111111111001011010100011111100001",
    "11111111110110110100011010101101101",
    "11111111110011010111001010111010100",
    "11111111101110010100000110110110100",
    "11111111101011110100100010000101100",
    "11111111110010011010101110110100101",
    "00000000000001101010001110010001010",
    "00000000010000011000100011011001000",
    "00000000010011110100111110001011001",
    "00000000001101110010110111001011111",
    "00000000000111000010001010011010010",
    "00000000000010110111000010001011010",
    "11111111111110011100100111101001001",
    "11111111111000001011001011010101011",
    "11111111110001011011010010001010111",
    "11111111101101011100110111111101101",
    "11111111101111001000111111010010110",
    "11111111110110000111011010010110111",
    "11111111111111100011011000001110011",
    "00000000000111110101111011111001100",
    "00000000001001111111011100001010001",
    "00000000000111100001110010111101000",
    "00000000000110010111101110011110001",
    "00000000000110101001000010011011101",
    "00000000000101110111001101110100001",
    "00000000000010110110111000111111000",
    "11111111111101101101010111110111101",
    "11111111111000110001001000101000101",
    "11111111110100101001110001111000101",
    "11111111110100000011000100001110001",
    "11111111111001100001010111110001011",
    "00000000000010001110011101101010001",
    "00000000001000001010000110000111101",
    "00000000001000001010100011011110101",
    "00000000000111011000011100100111001",
    "00000000001010001111101101100101000",
    "00000000001100101110100101001111000",
    "00000000001001011001001101110001011",
    "00000000000000011000001010101010100",
    "11111111111010000000011110110111111",
    "11111111111001000011001011111001111",
    "11111111111001101100001100010011010",
    "11111111111010010011101111100111110",
    "11111111111100010010000111100100000",
    "00000000000001110011100000111100110",
    "00000000000110111110111011010001101",
    "00000000000111011111001101001110111",
    "00000000000100001101001000101110110",
    "00000000000001000111100100000110101",
    "00000000000000111000010001010110011",
    "11111111111111010111111000111110100",
    "11111111111011010100010010110101001",
    "11111111110111011001011010000000111",
    "11111111110100101111110110000010101",
    "11111111110010111011110111010110001",
    "11111111110010011011010000101011011",
    "11111111111001001011010010111000000",
    "00000000001001011100101111011110100",
    "00000000011010110101110011111111110",
    "00000000100001101000100100111011001",
    "00000000011001000001111110011000010",
    "00000000001000001010110110111000010",
    "11111111111010111111000010001000111",
    "11111111110101110011000110001001011",
    "11111111110110111110001001111000111",
    "11111111111010010100010011011100100",
    "11111111111011100100100110110101110",
    "11111111111001110010001111010100001",
    "11111111111000011001001001011110100",
    "11111111111100011000011001011100101",
    "00000000000100100011110101100100111",
    "00000000001011100001100011010110001",
    "00000000001110110110111011101100110",
    "00000000001101000011111010111111000",
    "00000000000111100111100101111001001",
    "00000000000000101101101111110111000",
    "11111111111001110110010011100010011",
    "11111111110011110111100101011100110",
    "11111111101110100011001010011001100",
    "11111111101100111010001101111101001",
    "11111111110001001001000101001100001",
    "11111111111011001110110111000001110",
    "00000000000110100110001111101010100",
    "00000000001010011010001100000101100",
    "00000000000110111010111010111101000",
    "00000000000000010001000000110011010",
    "11111111111010110000000111111000110",
    "11111111111010101000011110111000010",
    "11111111111110000100010110101010001",
    "00000000000000111001110100010100011",
    "00000000000000111111110101101110011",
    "11111111111111110111011110010000000",
    "11111111111110011011111010001101010",
    "11111111111100110001111001101010111",
    "11111111111101101000000001110100101",
    "00000000000001001101101100111011101",
    "00000000000111010101111010110010100",
    "00000000001101010101010100111100011",
    "00000000001101111001010111011010111",
    "00000000001011000001001110100010111",
    "00000000000101110100000011100000000",
    "11111111111100011110000101101111110",
    "11111111110010101101010101011111111",
    "11111111101101101111011101111010011",
    "11111111110000010100010111101000000",
    "11111111111000011111100111111111011",
    "00000000000010001010001000111100001",
    "00000000001000101001101100110001010",
    "00000000001000111111000000011000101",
    "00000000000110010010011111111101010",
    "00000000000011011000101110001011111",
    "00000000000010110111001000100010101",
    "00000000000010100001100001011101110",
    "11111111111100011101101011011111110",
    "11111111110011111100111111101110110",
    "11111111101111011110111011100111001",
    "11111111110001011100010101000111110",
    "11111111110110010010000011011111011",
    "11111111111010011100011110011110011",
    "11111111111110000001100101100101100",
    "00000000000000000011110011011011011",
    "00000000000001100111100001101000000",
    "00000000000011101100010010101000011",
    "00000000000100110001111000001101011",
    "00000000000100001111010111100000000",
    "00000000000000111000001111001011010",
    "11111111111011011001110000000101111",
    "11111111110111101101010110110010101",
    "11111111110110100100011110001011111",
    "11111111110110100011001001100100001",
    "11111111111000110001010011010001110",
    "11111111111110110010010110011000010",
    "00000000000111001100010101110110100",
    "00000000001100100010001111111100100",
    "00000000001100101001101100101110010",
    "00000000000111001001110100111011110",
    "00000000000000101111000110011001011",
    "11111111111110010110110100000001000",
    "11111111111110110010010010101110010",
    "00000000000000100110110100000010100",
    "11111111111111100101111100110010001",
    "11111111111001011000011101011100000",
    "11111111110001000000011011010001110",
    "11111111101110011001101110001011110",
    "11111111111000001000010111001001001",
    "00000000001000010010101110101111011",
    "00000000010011101111100011111000010",
    "00000000010011000011000101010110010",
    "00000000001010001100110000010001111",
    "00000000000010011101100101011111110",
    "11111111111111111011001100101110001",
    "00000000000000010101110011111101111",
    "11111111111111000110101111010010101",
    "11111111111011100001011101110011010",
    "11111111110111110001011110110110001",
    "11111111110101101100110111101100100",
    "11111111110111010000110101010111101",
    "11111111111100111101001001000001101",
    "00000000000011011001110001000100011",
    "00000000001000101111111101011000010",
    "00000000001100100011011001111100100",
    "00000000001100111110010001010011011",
    "00000000001001101001000010011100100",
    "00000000000011000111011110010010001",
    "11111111111100010000010011010000011",
    "11111111110111001010111111111000110",
    "11111111110011110101100101000110111",
    "11111111110010000000001000011010000",
    "11111111110011100100111000010101000",
    "11111111111100100011011011001110000",
    "00000000001001010011010101100101000",
    "00000000010000001010111111111101101",
    "00000000001101000011000111111001101",
    "00000000000110100010111011101100111",
    "00000000000110000011111110110100001",
    "00000000001010011111101101000100100",
    "00000000001001100011001001110100011",
    "11111111111111001011110001001010000",
    "11111111110011010100000001001010100",
    "11111111110001111111111000101010010",
    "11111111111010101000100101111101001",
    "00000000000011101010100101100110100",
    "00000000000110110011100000011001111",
    "00000000000101110101000110111001001",
    "00000000000110011100000000101010100",
    "00000000001000011100011011110100011",
    "00000000000111011111011010101010110",
    "00000000000010101110001001101110010",
    "11111111111101011110111101011100011",
    "11111111111011111010110000010001110",
    "11111111111011101010011000100100000",
    "11111111111000111111100110100011000",
    "11111111110100111101111101110100011",
    "11111111110101100110010111011101000",
    "11111111111101011101010110010100100",
    "00000000000101000000100111010101010",
    "00000000000100110001010001100100101",
    "11111111111111111010011000110101101",
    "11111111111110000101100001011100000",
    "00000000000001111100010110010011111",
    "00000000000010110101101101110110100",
    "11111111111011010011001111000101100",
    "11111111110010011010101010001110111",
    "11111111101111101001101011110100010",
    "11111111110100111010011100100000101",
    "11111111111100011001100011010101100",
    "00000000000001010000011010011000100",
    "00000000000011111001011001001010000",
    "00000000000110101000101001111101010",
    "00000000001001101110010100001000000",
    "00000000001001001101000111010001111",
    "00000000000111000101001011111111110",
    "00000000000101011100101111010001000",
    "00000000000011010101001000100110101",
    "00000000000000101100111110100011111",
    "11111111111011110001111001111111010",
    "11111111110110000011000011100101001",
    "11111111110010111101101011001110110",
    "11111111110101111101000010111101010",
    "11111111111110101011111111110010000",
    "00000000001000111111101010001111101",
    "00000000001110100101001100111111110",
    "00000000001100011011000100001111110",
    "00000000001000000101011000111101110",
    "00000000000110111110010000001010000",
    "00000000000110100111010110000011010",
    "00000000000010001100111110010111001",
    "11111111111100000110110001001001010",
    "11111111111001101010111111111001001",
    "11111111111011011101011001100011001",
    "11111111111100100110100101100011011",
    "11111111111101000000101111000001001",
    "00000000000001000101100101011100000",
    "00000000000110011001110011001110100",
    "00000000001010100000001011010000110",
    "00000000001001110111010010000000110",
    "00000000000100010100101110110011011",
    "11111111111110111101101100001101011",
    "11111111111100010001000000000000111",
    "11111111111011100111100011010111010",
    "11111111111010101011000111111101010",
    "11111111111000101001110101011001001",
    "11111111110111000100001100110010000",
    "11111111111010001011111111011010101",
    "00000000000010001010010010011011111",
    "00000000001000111011011011011111100",
    "00000000001100110100110001011001111",
    "00000000001110010000001001110100010",
    "00000000001011001101110011010101101",
    "00000000000100100110111010011111011",
    "11111111111101010101100010011001000",
    "11111111111001100001100111111000111",
    "11111111111001101101010001110011001",
    "11111111111011110111100101111001100",
    "11111111111111010110010111011010010",
    "00000000000010010000010010001001100",
    "00000000000010101001111001011110101",
    "00000000000000110101001011000110011",
    "00000000000000011011011010110101110",
    "00000000000101100010010000010111100",
    "00000000001011111010101011101101011",
    "00000000001100011100010111100100011",
    "00000000000110111111000011111100111",
    "00000000000000000000101001010010001",
    "11111111111011100100110001011101111",
    "11111111111001011110000011010100001",
    "11111111110111100110001000100111111",
    "11111111110110010111101110010000001",
    "11111111110110101101011000001000011",
    "11111111111010011100000111011100110",
    "00000000000000000101001011101001010",
    "00000000000100111110110011000001000",
    "00000000000110111010011011000110101",
    "00000000000010101111010001000111000",
    "11111111111010000110111100011110011",
    "11111111110010010000101111001011111",
    "11111111110001011000100011001001001",
    "11111111110110110010010100011110001",
    "11111111111010100000011011001010011",
    "11111111111010001101101001011110010",
    "11111111111000110110101111010111101",
    "11111111111100001101010110011110111",
    "00000000000101000100010010001001111",
    "00000000001011111101001101101100001",
    "00000000001101011100011001111001000",
    "00000000001011100010101000010111101",
    "00000000001001000001101011011000101",
    "00000000000110000111111010011001101",
    "00000000000010110000011111100001001",
    "00000000000001011101111001000010110",
    "00000000000000011111111111011111110",
    "11111111111110110100011101001111001",
    "11111111111100101001111001101111001",
    "11111111111100001110101101001100011",
    "00000000000000110001110110111100101",
    "00000000000110111010110001110010111",
    "00000000001010100001111001111111100",
    "00000000001100000010010101001000110",
    "00000000001100011101001000100100101",
    "00000000001011000000111010010110000",
    "00000000000101000000101000111101000",
    "11111111111011001010110100100101111",
    "11111111110001100001001110111111011",
    "11111111101100010100010001010100111",
    "11111111101100001001001000010101100",
    "11111111101111110011011011011100010",
    "11111111111000111000001110000101010",
    "00000000000101010010110011010000110",
    "00000000001100101011101101100111101",
    "00000000001011010011111110001111010",
    "00000000000011101110110011100000000",
    "11111111111011011111111011000010111",
    "11111111110111111100110011001101101",
    "11111111111000000100101100100001000",
    "11111111111001011000110111000110001",
    "11111111111010101100100010100101101",
    "11111111111010100100001111010011001",
    "11111111111000000010000000100000101",
    "11111111110101111110100110000110100",
    "11111111111000100110000010010111110",
    "11111111111101110110110100011110111",
    "00000000000011110011010101011000101",
    "00000000001010000100100010101010110",
    "00000000001110001010011011011001010",
    "00000000001110011010101101001001001",
    "00000000001000001011110100000001100",
    "11111111111100110001010001111101000",
    "11111111110011011011001101010111011",
    "11111111110001110011110101010000100",
    "11111111110110101101010110111111000",
    "11111111111100000110000111001001011",
    "00000000000000100001101011101101010",
    "00000000000101000101001001000011000",
    "00000000001000001101001000010010001",
    "00000000001001000111000011010100001",
    "00000000000110100010001111110111111",
    "00000000000011100100010100101111001",
    "00000000000011000100001000110010000",
    "00000000000001001111100001101001000",
    "11111111111100000111110111100100101",
    "11111111110110100111100001100111001",
    "11111111110100110101110100111110001",
    "11111111111000100100100110110011010",
    "11111111111111001011011011000000101",
    "00000000000100111011000101010000011",
    "00000000000100100111010100011101110",
    "11111111111111100001000011000111011",
    "11111111111011000110100001101010110",
    "11111111111001100010111100011110010",
    "11111111111011101010000010001010101",
    "11111111111110001101110011101000000",
    "11111111111110101110011000001000111",
    "11111111111100111110111010011011010",
    "11111111111000100110111001001011111",
    "11111111110101110110111100010111111",
    "11111111110110110001000111001011000",
    "11111111111011000010100010101101011",
    "00000000000000011010001101010110011",
    "00000000000011111001001011001101001",
    "00000000000101101101000111001010011",
    "00000000000110101000111101101000110",
    "00000000000111000101111010010111011",
    "00000000000100101000010011100011100",
    "11111111111101011110000000010100000",
    "11111111110101110111111000011010000",
    "11111111110010000110011011100011101",
    "11111111110110010100001111001010111",
    "11111111111110101101000111101010001",
    "00000000000010111001010111011100110",
    "00000000000011011100110011100110100",
    "00000000000100010000011010011001100",
    "00000000000100111111001111101101111",
    "00000000000011110101111101100001010",
    "00000000000001000001110010001110110",
    "11111111111111010100000100101111010",
    "00000000000000110110101110111001111",
    "00000000000011000000100010100011011",
    "00000000000001100001000100110100110",
    "11111111111100010001010110100011010",
    "11111111111000010101001110000000011",
    "11111111111001011111101010000111110",
    "00000000000000100100000111010000011",
    "00000000001001111110000101001101010",
    "00000000001101110111110100111001111",
    "00000000001010011111111001101001011",
    "00000000000100111111111111001000100",
    "00000000000011101100010000100110100",
    "00000000001000110001000110000100010",
    "00000000001101110000011101110010000",
    "00000000001100101000011001000101101",
    "00000000000101100101000000110011010",
    "11111111111101101111011100110010001",
    "11111111111010100010001011111111011",
    "11111111111101001100111101000001100",
    "00000000000010100010110110101111101",
    "00000000000110101001011100010101101",
    "00000000001000000101001011111100001",
    "00000000000110101001101001001001110",
    "00000000000001110101100001101101001",
    "11111111111100110101001000001101001",
    "11111111111000100110101001000010111",
    "11111111110101011001110010111110101",
    "11111111110100001111101100001000010",
    "11111111110011001111000111110011001",
    "11111111110100011000000001111101111",
    "11111111111001010010010000111000000",
    "11111111111110111011100010001011110",
    "00000000000001010011101100010011110",
    "11111111111110111010010100111000111",
    "11111111111100010101001110011010100",
    "11111111111101000101010101001101010",
    "00000000000000010101011101110101110",
    "00000000000001111111011000110001011",
    "11111111111111100111111100101101101",
    "11111111111101100111001100001001100",
    "11111111111110010000111111000100011",
    "11111111111111000100000101011111100",
    "11111111111101010111011011011100110",
    "11111111111001111111011100000101001",
    "11111111111001111001101110011010101",
    "11111111111111100011100001001101110",
    "00000000001001010001100011100100001",
    "00000000010000011001001100000111000",
    "00000000001111101110011110110000010",
    "00000000001001001101111011001110111",
    "00000000000000101101001110000100100",
    "11111111111010000110111010111001110",
    "11111111110110000110100011001111110",
    "11111111110011100011100001101011100",
    "11111111110101010101011101110000010",
    "11111111111100100101101100010111100",
    "00000000000101011011001000110001100",
    "00000000001011001010101110011000110",
    "00000000001010111111001011111000110",
    "00000000000111010000010101111011000",
    "00000000000011011011001100001000001",
    "00000000000001100110000010111010100",
    "00000000000010010111001011011110110",
    "00000000000011101110101000001000110",
    "00000000000100000101101101100000001",
    "00000000000001111000010110010010101",
    "11111111111100100101111000001100111",
    "11111111110111010110101011101100001",
    "11111111110011101110111000101010101",
    "11111111110100010100011110100110011",
    "11111111111001111001101011111111000",
    "00000000000011010011101110110001100",
    "00000000001011110001010110110111111",
    "00000000001100100001001100111110001",
    "00000000000110100011110011101100111",
    "00000000000000110011101100110010000",
    "11111111111111110010111100010011111",
    "00000000000001110001011001111101010",
    "11111111111111101011101001100011101",
    "11111111111001111111110010001000010",
    "11111111110110010011111101001101001",
    "11111111111010100111001010011100110",
    "00000000000100001011001001000110001",
    "00000000001010101010000101001000000",
    "00000000001011010011001100100000000",
    "00000000000110101001110010110111010",
    "00000000000001000100000111100111111",
    "11111111111110101111010101100110000",
    "11111111111101101000001111000001000",
    "11111111111011110001010100100011011",
    "11111111111010010010100001001010000",
    "11111111111011111011001100111000111",
    "11111111111111101011101001011100111",
    "00000000000001100101001010111010100",
    "11111111111111101011100100001011100",
    "11111111111011110111000100011111110",
    "11111111111100011011101110011011100",
    "00000000000001011001000110010010101",
    "00000000000011110011010111011101100",
    "00000000000000110000001011101110110",
    "11111111111011011100011010010101110",
    "11111111111000010000010000011001000",
    "11111111111000100001101101111111001",
    "11111111111001001000110010000111011",
    "11111111111000001100110001001101111",
    "11111111110111000000111000101110100",
    "11111111111000110111100101111011011",
    "11111111111101001110111111000010110",
    "00000000000001101101100000000011111",
    "00000000000101010100011011011100000",
    "00000000001000110000111011101000111",
    "00000000001011001001101101001011000",
    "00000000001100000101100101101010010",
    "00000000000111111011011100010000101",
    "11111111111110111011111100100001001",
    "11111111110110010001110101001111011",
    "11111111110010111110010111111111001",
    "11111111110101111111011101011101110",
    "11111111111011111000111100111011111",
    "00000000000010101110111110010111111",
    "00000000001001000010010110011001011",
    "00000000001110001010100010100000101",
    "00000000010001000111000010001001010",
    "00000000001101100011100010101010010",
    "00000000000101010010010100001000010",
    "11111111111011100101010001011110011",
    "11111111110101101010000110010111110",
    "11111111110110010010001100001111010",
    "11111111110111110011111110000100000",
    "11111111111000110011101111111010011",
    "11111111111010110110111100101001110",
    "00000000000000100101001101110001100",
    "00000000001001110100011111111000001",
    "00000000010000110011111110010101001",
    "00000000010001111001000110111111110",
    "00000000001100111100100011000110100",
    "00000000000101011111000111100011111",
    "00000000000000010000100111101000011",
    "11111111111101100101001000001011011",
    "11111111111100011001010011000000010",
    "11111111111010111000110010000111000",
    "11111111111011010110000101101100101",
    "11111111111110001001001101011001001",
    "00000000000000001110110001010000111",
    "00000000000001001111100110001110111",
    "00000000000010011100111001100011011",
    "00000000000111011000011010001101100",
    "00000000001110001101110111000000110",
    "00000000001111000001101000101110001",
    "00000000001001111010011110001000100",
    "00000000000001110111011110010100111",
    "11111111111100000111101000101101101",
    "11111111111011000100010011010000011",
    "11111111111011010001000101111110101",
    "11111111111010100111110011000000100",
    "11111111111011101110000010101001001",
    "00000000000000101110001111101110110",
    "00000000000110011110011110011000101",
    "00000000001001100001101001110100111",
    "00000000001000010001101011000010001",
    "00000000000010010011011111010010110",
    "11111111111101111101110101101100100",
    "11111111111111101100100000111100110",
    "00000000000100001111101010011011000",
    "00000000000101101000101110001100111",
    "00000000000000100111001110010001111",
    "11111111111000111001100111000010011",
    "11111111110101111101010000010100111",
    "11111111111001110111111000000101111",
    "00000000000001010010011101001100100",
    "00000000000111101001000010100000000",
    "00000000001010001110010011001111011",
    "00000000000111110011010010010100001",
    "00000000000010011110010100000011110",
    "00000000000001001101010011111101000",
    "00000000000100111100100111000001110",
    "00000000000110001010100101011111100",
    "00000000000000111101100100100101001",
    "11111111110111111101111110011001111",
    "11111111110010110101100001100110101",
    "11111111110111001111010001010011011",
    "00000000000010110101010000010100000",
    "00000000001101111000111001100010000",
    "00000000010010000000010011000000010",
    "00000000001111101000101100001110010",
    "00000000001010010101101101011011111",
    "00000000000110011001011101011000111",
    "00000000000101001011000010110010110",
    "00000000000100010010101101000001100",
    "00000000000011001011110110110000010",
    "00000000000000001001011101111001110",
    "11111111111100111001001100111110101",
    "11111111111100101010000000011111111",
    "11111111111101110110111101100001101",
    "00000000000001101010000100110010000",
    "00000000000110111001100110000001011",
    "00000000001011001111110011100001010",
    "00000000001101101110111010111110011",
    "00000000001100111101011010010100101",
    "00000000001011110111000010101110111",
    "00000000001010000111001000011101101",
    "00000000000011101101111111001110100",
    "11111111110111111110001000111011000",
    "11111111101101010100100000010110011",
    "11111111101101100100101101001101000",
    "11111111111000011101101010101110011",
    "00000000000110100000010011000111001",
    "00000000010000010111001011001010000",
    "00000000010001011011100010100111101",
    "00000000001100011000100000110101001",
    "00000000000111000111100000010100011",
    "00000000000101000011001110001011100",
    "00000000000011101001011100001001001",
    "11111111111110110110110000011010110",
    "11111111111000101111111010001000000",
    "11111111110101010001100001000110010",
    "11111111110110111100001000101001011",
    "11111111111010111111010000000010111",
    "11111111111011110000111100010010000",
    "11111111111011000010100001101111000",
    "11111111111010100010011001100001011",
    "11111111111100110111000111100001111",
    "00000000000010010110011101011110110",
    "00000000000101101010101111110000001",
    "00000000000010011001010001011001110",
    "11111111111010110010011110011011011",
    "11111111110101011010110011100010101",
    "11111111110110000110000100000111000",
    "11111111111010001001001110010101011",
    "11111111111111010010101001011110010",
    "00000000000010010011010100110110011",
    "00000000000010101101011000001101111",
    "00000000000100111001011010110100101",
    "00000000001001010001000111010100100",
    "00000000001100010101101000011101010",
    "00000000001010001011000001010101110",
    "00000000000011001000011010001000100",
    "11111111111100011101000000011100110",
    "11111111111000100100001100110111111",
    "11111111110111100110001101000110110",
    "11111111110111000101001010110000011",
    "11111111111001000010000101111101110",
    "11111111111100111010000001011101010",
    "11111111111110010111001010100111101",
    "11111111111111000010001101010100110",
    "00000000000000010000001101101101110",
    "00000000000010001010010110101111100",
    "00000000000011001101101011011001110",
    "00000000000001110111010100001010000",
    "00000000000000010010010100001011110",
    "11111111111111011001110010111111110",
    "11111111111111101001000111111001000",
    "00000000000000011100010101010010111",
    "11111111111111011011100100000011011",
    "11111111111011100111010100110001010",
    "11111111110111010010000110000111001",
    "11111111111001001110101011110101100",
    "00000000000011010100010111011100111",
    "00000000001110010001011011100010100",
    "00000000010001000010110011001011100",
    "00000000001001101000000111100011001",
    "00000000000000110111000000000011011",
    "11111111111101001001110111110010001",
    "11111111111100011101111111011001011",
    "11111111111001101110011110111001110",
    "11111111110011100110111000110100111",
    "11111111101110101101101000111110000",
    "11111111110001101011001011111000001",
    "11111111111010100110011111010011101",
    "00000000000011011001011101100110110",
    "00000000001000010110101111011001010",
    "00000000001001010111011011101101101",
    "00000000001000111011011111100001100",
    "00000000001001000001000010111001010",
    "00000000001000011001110110011111010",
    "00000000000101011001011101111000110",
    "00000000000000111010011001110011000",
    "11111111111100001110101011100111101",
    "11111111110101111100101010001100010",
    "11111111110010100001010110010001100",
    "11111111110011111110100111011111111",
    "11111111111001001101101110010100100",
    "00000000000000011100011110101000001",
    "00000000000101110111111000110001110",
    "00000000001001011100001111001101001",
    "00000000001010110101000101110000001",
    "00000000001000010011101111111011011",
    "00000000000010110011010011001000100",
    "11111111111101110110111100111100000",
    "11111111111100011000011110111001110",
    "11111111111010101101000101011101001",
    "11111111110111110010100000000101001",
    "11111111110111100011001001100100001",
    "11111111111101011101010000111000101",
    "00000000000110101111101111011010100",
    "00000000001001111101001011011111000",
    "00000000000100111001110110101111101",
    "11111111111110111000100010100111100",
    "11111111111111000010110010100001011",
    "00000000000010111001010111110101011",
    "00000000000011110100001101101001000",
    "00000000000000101010101000010100010",
    "11111111111110001011010000000001010",
    "11111111111110100110100010111011001",
    "11111111111111000111110010011110101",
    "11111111111100100100010100101001010",
    "11111111111010001000011100011111011",
    "11111111111110101110101011110011111",
    "00000000001001100101010001000000010",
    "00000000010001010111101100111011110",
    "00000000001111000111011110011101010",
    "00000000000110101100010110110101001",
    "00000000000000111111110111110011111",
    "11111111111110101101101110101011110",
    "11111111111010111110111001101100000",
    "11111111110100001000101000001101000",
    "11111111110000101101110011011010000",
    "11111111110110011100000001011100101",
    "00000000000000010011011010111110000",
    "00000000000110101001110001111000001",
    "00000000000111101100010100010000000",
    "00000000000111010000110000010111110",
    "00000000001000101000010010110000110",
    "00000000001001011011010110011111100",
    "00000000000111010010100101111000100",
    "00000000000001001010111101101011010",
    "11111111111001000111100010111010001",
    "11111111110011110100111111111111111",
    "11111111110100110101000111000011111",
    "11111111111101010111100000000111110",
    "00000000000111100100110000010111010",
    "00000000001100010011000100111111101",
    "00000000001010001111010101001100010",
    "00000000000101011000110000110011100",
    "00000000000011001001010110110110110",
    "00000000000010000011111101011001100",
    "00000000000000001100001101101101111",
    "11111111111101001111100010011101111",
    "11111111111001100101111110100110110",
    "11111111110110111011000110100010111",
    "11111111110110110011101001111001010",
    "11111111111010001010110000111110100",
    "11111111111110011010010110000011001",
    "00000000000001110010011100100110001",
    "00000000000110000111000000001011010",
    "00000000001010010010101101110101000",
    "00000000001110001101101110010100001",
    "00000000001111011110110011110001111",
    "00000000001001110011011101000011111",
    "00000000000001001111000010100001000",
    "11111111111100001001011010111010000",
    "11111111111100001010000101011011011",
    "11111111111100111010110101101000111",
    "11111111111010101001010011011001101",
    "11111111110110101100000110010011110",
    "11111111110100011110101101100000001",
    "11111111110110111100011011000011101",
    "11111111111011011100110101011100111",
    "00000000000000101001000011101010001",
    "00000000000111001110001011101100001",
    "00000000001100000001110101101001111",
    "00000000001011011010100000010110010",
    "00000000000110010001110111111011110",
    "11111111111110100101111011101011101",
    "11111111110110110110011000001101110",
    "11111111110010000101101111100110010",
    "11111111110010111110001100001011000",
    "11111111111000010110001010100110100",
    "11111111111101010110110100011110010",
    "00000000000010011010101110110101110",
    "00000000000111110111101101001111011",
    "00000000001010111011110001111001011",
    "00000000000111011100111110111011100",
    "11111111111101001101100111110101101",
    "11111111110101111111101110011000000",
    "11111111110101111011010101100001101",
    "11111111111010000001100001110010010",
    "11111111111101010101010010111111001",
    "11111111111101100010100000101010101",
    "11111111111100101001100101000011100",
    "11111111111001101011010111110001001",
    "11111111110110101100000111011111001",
    "11111111111000110101000101101101010",
    "00000000000000010101100010001100100",
    "00000000000111001101000101101000111",
    "00000000000110001011101000010001011",
    "11111111111111111001111101111110101",
    "11111111111011100101100111001001010",
    "11111111111011010100011111100101000",
    "11111111111101001001000001001101011",
    "11111111111101100010010100000001101",
    "11111111111100001100010000000000011",
    "11111111111011000010010001111110100",
    "11111111111011110101110110100011111",
    "11111111111111010001110001111011101",
    "00000000000001011110101010000101111",
    "00000000000001000101001000001011010",
    "00000000000001111000011000000111100",
    "00000000000100100110000111000100111",
    "00000000000110000111010001001000000",
    "00000000000010001101110100010100000",
    "11111111111010000010110110000111100",
    "11111111110100011111010100001010101",
    "11111111110100110000011011000001111",
    "11111111111001011110000001101100001",
    "11111111111101001110111101010001011",
    "11111111111111001010010011100000100",
    "00000000000001110100000010110010010",
    "00000000000101110010011101011000010",
    "00000000001010110101010110111001110",
    "00000000001101011111011011110001100",
    "00000000001011000011101010111101100",
    "00000000000100011101111101110000110",
    "11111111111101010111111011011000110",
    "11111111111010100000101100100000111",
    "11111111111001101110001011000100010",
    "11111111111001100011100111101110011",
    "11111111111011000101010100110101001",
    "11111111111110101011110110010011101",
    "00000000000100001000001001001010010",
    "00000000000111111001111001111100111",
    "00000000000111111001100100110000110",
    "00000000000110111010110001010110111",
    "00000000000110011011001001000100100",
    "00000000000110011011011001001101101",
    "00000000000100011010010101111100000",
    "00000000000000110000100101111100110",
    "11111111111011100001001010101010011",
    "11111111110100000011110010001010100",
    "11111111101111001111100101000000111",
    "11111111110011001000100011110010101",
    "11111111111111010110001010111001011",
    "00000000001011001001110111010010111",
    "00000000001110010100011010101110110",
    "00000000001011010111011010110011001",
    "00000000000111101010101001000100100",
    "00000000000111101110000100011011011",
    "00000000001001011000010100110101011",
    "00000000000110100001110101101001000",
    "11111111111101111101101111110010101",
    "11111111110011010011011000011101011",
    "11111111101101100100011101010101100",
    "11111111101111011110000000111110111",
    "11111111110110111100111111010100000",
    "11111111111111110100101110011100011",
    "00000000000101001101000010110011101",
    "00000000000110110000101011010111010",
    "00000000000101001011111001101010111",
    "00000000000000110000011001100001111",
    "11111111111101011100010000101011111",
    "11111111111100010100010000100101110",
    "11111111111010010111000010110101100",
    "11111111110110001001100111111010111",
    "11111111110011100001100101110101110",
    "11111111110100101101000010000111011",
    "11111111111001010000110111000110110",
    "11111111111110111001101101110111110",
    "00000000000011001100110100011000011",
    "00000000000101101000101110010000111",
    "00000000001001101010101111101001110",
    "00000000001101101010001110110110011",
    "00000000001101101001110000100010111",
    "00000000001001000101010100011110100",
    "00000000000000100011111110111000010",
    "11111111111000000101110100100101011",
    "11111111110100100100101000100011001",
    "11111111110101101010010110110001110",
    "11111111111000001001000111001011011",
    "11111111111011011110100010111101101",
    "00000000000010010011000101110110000",
    "00000000001010110111110110011001011",
    "00000000010001010010100010111101110",
    "00000000010001011000000110111000011",
    "00000000001001111011011001010110101",
    "00000000000001101000110011000110010",
    "11111111111101100110010110010100110",
    "11111111111011001001100011001101011",
    "11111111110111000110001101011101100",
    "11111111110001111101110001011110100",
    "11111111110000001001001111111100101",
    "11111111110100001111101110101111001",
    "11111111111100000100100101101011110",
    "00000000000100110011010011010000101",
    "00000000001011011110100000000100011",
    "00000000001101101100000010010111110",
    "00000000001000110010110100001011100",
    "00000000000000110101001010110001101",
    "11111111111011101110001100110000000",
    "11111111111010001010001000100000010",
    "11111111111010101101000100010110100",
    "11111111111010001101111011110000011",
    "11111111111001011110000111001011010",
    "11111111111010101101000111100000100",
    "11111111111110000111101001110000100",
    "00000000000101000101101011001010001",
    "00000000001011101000010110010011111",
    "00000000001100110011011010000110000",
    "00000000001000000100010110111110111",
    "00000000000010100111110101011001100",
    "00000000000000100010111111111000110",
    "00000000000000101000100110110111000",
    "00000000000000010001100110000010000",
    "11111111111101010100011110100001101",
    "11111111111001001111110101100000100",
    "11111111110110100101000011110100110",
    "11111111110110011000010111111010100",
    "11111111111010100011101100010010110",
    "00000000000001110110000001000000100",
    "00000000000111000001010101111100010",
    "00000000001001000101100110100010010",
    "00000000001010010100101000001110000",
    "00000000001010011110100110111010010",
    "00000000001000001111010000010110010",
    "00000000000001100100100101111111110",
    "11111111110111001101011001010101001",
    "11111111101111110110000010110100000",
    "11111111110001100001011011011111101",
    "11111111111001100001111111110100101",
    "11111111111111100000100011000010110",
    "00000000000010001111011100111001001",
    "00000000000010110001010111110101100",
    "00000000000100011110100101100110101",
    "00000000000111001001100110100101010",
    "00000000000110110001011011001001011",
    "00000000000010000011011100001000110",
    "11111111111010101010111100111001111",
    "11111111110101000001010110001011100",
    "11111111110100000000111001011101001",
    "11111111110110001111100101011111010",
    "11111111111001010001001001011000010",
    "11111111111011011101101000100010011",
    "11111111111111000010001001101010001",
    "00000000000101011010101100100110111",
    "00000000001100000101000110001010110",
    "00000000001110110001010111001101111",
    "00000000001100000111000010001101101",
    "00000000000101110000011001010010010",
    "11111111111111100001001111100011001",
    "11111111111100001101001101011110011",
    "11111111111011110000010010101101000",
    "11111111111001111101100110101110010",
    "11111111110110110110010110100100100",
    "11111111110111100010100011001101001",
    "11111111111011110101011100110100001",
    "00000000000001011011110000010101001",
    "00000000000101100111010110000011010",
    "00000000001000010011110110111100101",
    "00000000001010101111011101000110001",
    "00000000001001001001100101001011111",
    "00000000000010001100110101011000110",
    "11111111111001011000111010111101001",
    "11111111110101010100101000111101100",
    "11111111110101100000010001111000011",
    "11111111110101011100110111000110010",
    "11111111110111001010110100001101110",
    "11111111111010101111001001010011100",
    "11111111111111100000010011001000110",
    "00000000000011110010100101010000101",
    "00000000000101011111011100001010011",
    "00000000000111001100111010100111110",
    "00000000001001111001011100001000011",
    "00000000001000101011000101000101000",
    "00000000000000000111000010010110110",
    "11111111110101100110111110101111110",
    "11111111110000000101111110011101000",
    "11111111110000111101100001000101100",
    "11111111110101010010110101010010111",
    "11111111111000110110111011110101000",
    "11111111111011111101100011001100010",
    "00000000000000110111011101110000010",
    "00000000000101000110111001110100100",
    "00000000000110011011110010111110011",
    "00000000001000001111010100010011010",
    "00000000001010101001000000011101010",
    "00000000001010011010111001100100011",
    "00000000000011110110110001100111010",
    "11111111111001101001001111111000010",
    "11111111110100100001001000101001000",
    "11111111110110111110000110110001101",
    "11111111111100011111100011100010010",
    "11111111111110110000011000101100000",
    "11111111111111000110100010010010000",
    "00000000000011111101110111101010010",
    "00000000001100100011111011101010110",
    "00000000010010100100010001000001001",
    "00000000010000100010010110001011001",
    "00000000001000011101110111100111110",
    "00000000000000011110110010001111011",
    "11111111111011010010110000100111000",
    "11111111111001100011001010010000011",
    "11111111111001101011101101011001001",
    "11111111111011001111011010110001101",
    "00000000000000010100010101000001000",
    "00000000000111010110011011111101011",
    "00000000001011101011101011110010100",
    "00000000001001100110011100100100100",
    "00000000000001111111111011010001011",
    "11111111111010111000000101111000001",
    "11111111111000001001100010011110110",
    "11111111111001100101011101000101100",
    "11111111111011010010101011010111100",
    "11111111111100000001111101001110110",
    "11111111111011000101100111001101110",
    "11111111110111011011110111010101000",
    "11111111110110001001000100011111010",
    "11111111111000110011010000010101101",
    "11111111111100100101011000110011110",
    "11111111111111111101001111001010001",
    "00000000000001111000000111100100000",
    "00000000000100011110100101010110110",
    "00000000000111100010111110101111100",
    "00000000001000001100111001110101100",
    "00000000000101000000001110110001001",
    "11111111111111101110001000011110111",
    "11111111111011110000110010111101010",
    "11111111111000110110011101100010101",
    "11111111110110101010101100011101000",
    "11111111110101110001111111110011000",
    "11111111110111010011011001010101010",
    "11111111111101110000100010001110111",
    "00000000000101011101100100000100011",
    "00000000001001101001000000001010110",
    "00000000001001011010001110100100000",
    "00000000000111000010010001101101001",
    "00000000000101011001001010011101001",
    "00000000000011001011101101001001001",
    "11111111111111100101001000010101111",
    "11111111111011100000000001010111010",
    "11111111110111101000100101110011001",
    "11111111110100001111011000101011111",
    "11111111110011000011101100110010011",
    "11111111110111001010000100101000101",
    "00000000000000010100001111011000100",
    "00000000001001000001100001111000010",
    "00000000001101011111100111000111001",
    "00000000001110111001001001011110101",
    "00000000001110111001000110000110000",
    "00000000001011010001000111010101101",
    "00000000000001111000011010110010000",
    "11111111110111100000001110011000110",
    "11111111110100000101001111101011110",
    "11111111111010001101100110100000111",
    "00000000000010110010101001000101011"
  );

  constant PKG_OUTPUTSAMPLESFI_CONCAT : std_logic_vector(87219 downto 0) := (
    "11111111110111101001100100111110010" & 
    "11111111110010001100111000111011001" & 
    "11111111110100111110011101011000110" & 
    "00000000000000101001010000011001011" & 
    "00000000001011111110100111000111111" & 
    "00000000001111100000100111000100110" & 
    "00000000001110011101010001011011010" & 
    "00000000001101110100010111100010000" & 
    "00000000001110101111100111101101110" & 
    "00000000001100010000100001101110101" & 
    "00000000000101100000101001000011010" & 
    "00000000000001000001110110101011111" & 
    "00000000000000101111010000010000111" & 
    "00000000000011001010111100001111101" & 
    "00000000000100100010001001101100110" & 
    "00000000000000100000001111001100100" & 
    "11111111111011000010001101110010010" & 
    "11111111111010111001101110010111010" & 
    "00000000000010010000100010001110110" & 
    "00000000001011110000101010110111111" & 
    "00000000010000111110000001000100100" & 
    "00000000010000001110100111111001100" & 
    "00000000001010111100101101101011111" & 
    "00000000000101001100110110110111001" & 
    "00000000000000000101110110011001000" & 
    "11111111111011110010011100110011001" & 
    "11111111111000101010001101010011000" & 
    "11111111110011010000011100111001111" & 
    "11111111101101110001011101010011101" & 
    "11111111101101111111010001111110011" & 
    "11111111110101100010001101010001011" & 
    "00000000000001011110100010110001010" & 
    "00000000001010001100010101100011001" & 
    "00000000001100001000111100111011010" & 
    "00000000000111100010100001001110010" & 
    "00000000000001110000000011001110000" & 
    "11111111111111000010000010100000011" & 
    "11111111111101010010011011011101100" & 
    "11111111111011110100110111110111000" & 
    "11111111111000001111110110010101001" & 
    "11111111110100100000111011011100011" & 
    "11111111110101110001000010010010010" & 
    "11111111111100101001010000111011001" & 
    "00000000000110011110011001000101001" & 
    "00000000001100111111101101111111000" & 
    "00000000001101100011000000101111100" & 
    "00000000001000111111010110111111001" & 
    "00000000000000111111100111100111010" & 
    "11111111111011101101101100100001000" & 
    "11111111111010111110001110101101100" & 
    "11111111111100011000110110100010010" & 
    "11111111111100011011101100100001111" & 
    "11111111111010010011011011011100001" & 
    "11111111111001011011000010100000101" & 
    "11111111111011001111001010011001100" & 
    "11111111111110000101010000010000000" & 
    "00000000000000110011100110000101110" & 
    "00000000000101001010110101010011100" & 
    "00000000001101010100011011011011011" & 
    "00000000010010110001111001001011010" & 
    "00000000001111010001010010100010000" & 
    "00000000000010101001101000010101010" & 
    "11111111110101110000010001100110101" & 
    "11111111110001101001101110111110001" & 
    "11111111110110000110111110010010001" & 
    "11111111111011111001001000000100100" & 
    "11111111111110111000101000010101011" & 
    "00000000000000100111111001001110100" & 
    "00000000000011101101011111101111110" & 
    "00000000000100111110101111100101111" & 
    "00000000000010010011000111000111000" & 
    "11111111111111010000110011000001000" & 
    "11111111111110110111101000110001100" & 
    "00000000000000100110100010010000000" & 
    "00000000000001100111001010010110100" & 
    "11111111111111101101111011101010011" & 
    "11111111111101111101001100110001000" & 
    "11111111111101001011010010100001110" & 
    "11111111111101000100001010111001101" & 
    "11111111111101110101011100101001111" & 
    "00000000000000111110011010001010100" & 
    "00000000000110000101100001100100101" & 
    "00000000001010000000011010110100110" & 
    "00000000001010010100101100000111001" & 
    "00000000000101000001011010001110000" & 
    "11111111111101011011110110000011100" & 
    "11111111111011001110100110111001001" & 
    "11111111111110101011010000001110100" & 
    "00000000000011001100101110111101010" & 
    "00000000000011010010010101110100010" & 
    "11111111111110000100011010111011100" & 
    "11111111111000110111000001000101010" & 
    "11111111110101111001101000000100000" & 
    "11111111110110111101000001100110110" & 
    "11111111111011000011101001101110001" & 
    "00000000000000111011010111110101100" & 
    "00000000000110001110101111100011111" & 
    "00000000000110101010101111111011111" & 
    "00000000000011100001011111110111011" & 
    "11111111111110100011010001001011011" & 
    "11111111111001110000010001010010100" & 
    "11111111111000100000101010111010100" & 
    "11111111111011110100100011001010111" & 
    "00000000000001010001110010111101000" & 
    "00000000000001000000101011101010001" & 
    "11111111111100001000110110101111001" & 
    "11111111111010000111111000110010010" & 
    "11111111111110101100001100001100010" & 
    "00000000000110010101010001011010101" & 
    "00000000001011011001001000111011001" & 
    "00000000001011011000111111101101101" & 
    "00000000000111101001101111001110101" & 
    "11111111111110101000010000110100000" & 
    "11111111110100000010011101001111110" & 
    "11111111110000010010001110110000101" & 
    "11111111110111111110101100000010001" & 
    "00000000000100001101100101101011001" & 
    "00000000001001110010011001001010111" & 
    "00000000000110100010111011100101001" & 
    "00000000000001110001000100001101001" & 
    "00000000000001111111101010000101111" & 
    "00000000000111111000100110110110101" & 
    "00000000001011011100010001111101111" & 
    "00000000001000001100111110010110110" & 
    "11111111111111001101100111110100101" & 
    "11111111110101101010111100100101001" & 
    "11111111101111101000100100101101110" & 
    "11111111101110011110000111111001010" & 
    "11111111110011010100101100100110100" & 
    "11111111111010000110111101100010101" & 
    "11111111111110110110000000111100110" & 
    "00000000000010011010111101001011010" & 
    "00000000000101011000000110110101001" & 
    "00000000001001011000000110100000100" & 
    "00000000001011101100001010110101010" & 
    "00000000001000100010111110011100010" & 
    "00000000000001001001100010111111011" & 
    "11111111111001000100001001000011000" & 
    "11111111110011111001110101110011111" & 
    "11111111110001000101011010000010010" & 
    "11111111110001001100101010101001001" & 
    "11111111110010011100001010110101000" & 
    "11111111110011001010010100100101010" & 
    "11111111110111010010100010111110101" & 
    "11111111111111011111111110100101110" & 
    "00000000001000010100101010001000000" & 
    "00000000001100100110011101100111110" & 
    "00000000001001100100011010111001011" & 
    "00000000000100000010000000010010010" & 
    "11111111111111010010000010110100010" & 
    "11111111111100000110000001111011100" & 
    "11111111111010001010001001101010101" & 
    "11111111111001010101110010101010111" & 
    "11111111111010001110111000110001110" & 
    "11111111111011110000000101100100010" & 
    "11111111111011010110001110101001000" & 
    "11111111111010101110000000101010101" & 
    "11111111111111001111111001110000110" & 
    "00000000001010001110100010100110010" & 
    "00000000010011101000110001111010011" & 
    "00000000010010110011011110000000011" & 
    "00000000000110100000111111111100111" & 
    "11111111111000011101111110011101011" & 
    "11111111110100010111000111011001100" & 
    "11111111110110111111010100001001010" & 
    "11111111110110000000111101110100111" & 
    "11111111110000100111110111111010100" & 
    "11111111101110000101001010011111010" & 
    "11111111110101100100010100111001001" & 
    "00000000000010101000111110011100110" & 
    "00000000001011111111001011001110000" & 
    "00000000001101000000101010101101110" & 
    "00000000001001000010010001001000110" & 
    "00000000000100101111010101100000000" & 
    "00000000000000010111000011011101101" & 
    "11111111111011100100001101110010101" & 
    "11111111110110111010011001110011100" & 
    "11111111110011001011111010011001011" & 
    "11111111110100100001001001000100011" & 
    "11111111111010000011101010011010010" & 
    "00000000000000000111111010101100110" & 
    "00000000000101011000011010011011000" & 
    "00000000001001011000011101001001110" & 
    "00000000001100000111001111111110010" & 
    "00000000001100010000000100010000100" & 
    "00000000001000000100001110000110001" & 
    "00000000000001010001100011111111010" & 
    "11111111111010111100110100111000010" & 
    "11111111110111100001100101011000111" & 
    "11111111110110110100101111100111000" & 
    "11111111111010010100011100011100000" & 
    "00000000000000010000001010011110101" & 
    "00000000000100001110100000101000010" & 
    "00000000000110011111101101000000010" & 
    "00000000000111001110010010111111100" & 
    "00000000000111001101111110100110000" & 
    "00000000000111100010111110011101101" & 
    "00000000000110110101100010010110101" & 
    "00000000000101100100100011110100001" & 
    "00000000000011111000100110000001001" & 
    "00000000000000100101001011000011101" & 
    "11111111111011100100110010110111100" & 
    "11111111110110111010101110110101100" & 
    "11111111110100100111010010010010111" & 
    "11111111110110001001011111101010001" & 
    "11111111111100110110011111110110110" & 
    "00000000000101001111010001011100110" & 
    "00000000001001100111000010101001011" & 
    "00000000001000100111100001110111100" & 
    "00000000000011101101100100101001100" & 
    "11111111111101110011000000001000010" & 
    "11111111111011000101011101011010000" & 
    "11111111111011110100010011111111100" & 
    "11111111111100101110010111010111100" & 
    "11111111111010110011110000001011011" & 
    "11111111111000010110111101111011100" & 
    "11111111111011011000000001100100110" & 
    "00000000000010001100101010111001000" & 
    "00000000000110100111011110000001000" & 
    "00000000000100100011010101110010110" & 
    "00000000000000101010000110101001001" & 
    "00000000000001101000110101100111101" & 
    "00000000000100101101100101000110011" & 
    "00000000000101111001011101001101110" & 
    "00000000000011101100010100110001101" & 
    "11111111111110110000011000001011001" & 
    "11111111111000011010111010011001001" & 
    "11111111110010000011000000101111000" & 
    "11111111101111110110011101000110011" & 
    "11111111110100011101110110001111000" & 
    "11111111111100000101101001010000101" & 
    "11111111111111010010001000101111000" & 
    "11111111111110000011000110100110011" & 
    "11111111111110010010001101101010000" & 
    "00000000000001100010100000111110100" & 
    "00000000000101011111110010010110100" & 
    "00000000000110001100101111111100011" & 
    "00000000000010100100101101100111010" & 
    "11111111111101111011011100010000100" & 
    "11111111111000010110011110000111100" & 
    "11111111110011000101101000011000010" & 
    "11111111110100001010111000110000111" & 
    "11111111111100010111010100110110001" & 
    "00000000000101101001000110000011010" & 
    "00000000001001011000101011110110100" & 
    "00000000000111010010110100001110100" & 
    "00000000000101010111101101110010000" & 
    "00000000000101111011111111001000000" & 
    "00000000000101000000011010000000010" & 
    "00000000000001101110101100100101000" & 
    "11111111111101011001010000110110011" & 
    "11111111111001110001000110010100001" & 
    "11111111111000001001100111001111100" & 
    "11111111111010111110011101110101001" & 
    "00000000000000101010100100110110110" & 
    "00000000000100101000110001010100001" & 
    "00000000000100010010011100000101001" & 
    "00000000000001101000110111011010101" & 
    "00000000000001111110000011011011100" & 
    "00000000000100101100101110001000001" & 
    "00000000000100000100011110101100011" & 
    "11111111111111001101101101000110010" & 
    "11111111111000111110000010001010100" & 
    "11111111110110010110101011000111110" & 
    "11111111110111000010001111101001010" & 
    "11111111111010100111011011001111101" & 
    "11111111111111111011011001011110101" & 
    "00000000000011111111000000111000001" & 
    "00000000000110001000000110011110011" & 
    "00000000000101100001000111100000010" & 
    "00000000000010110111110101101001010" & 
    "00000000000001111100101100100111111" & 
    "00000000000010100111010010011111101" & 
    "00000000000011010101011000111100010" & 
    "00000000000010011100001101000000000" & 
    "11111111111111100100111110111111111" & 
    "11111111111100100111101001110001100" & 
    "11111111111100000100100111011000011" & 
    "11111111111110111100101100000111100" & 
    "00000000000010100110011010010001101" & 
    "00000000000100000100110111111101011" & 
    "00000000000100000000011010001101100" & 
    "00000000000100000010001101000100000" & 
    "00000000000110011001000111001100111" & 
    "00000000000110101100000101001011010" & 
    "00000000000001011101010010101011100" & 
    "11111111111011010010100110101101100" & 
    "11111111111001010000101101101010001" & 
    "11111111111100111100101001001001111" & 
    "11111111111110011000111100110101010" & 
    "11111111111010010101101010000111110" & 
    "11111111110110001001101110111011101" & 
    "11111111110100001101101101101010001" & 
    "11111111110101101111111101110010011" & 
    "11111111111000000000100001111000000" & 
    "11111111111011000111111001010100000" & 
    "11111111111111111100000101001001110" & 
    "00000000000101011001100111010010101" & 
    "00000000001000100000000100001011100" & 
    "00000000000101110010001001100111100" & 
    "11111111111111101110110101101010110" & 
    "11111111111001110101011100110111001" & 
    "11111111110111000010110100101111111" & 
    "11111111111010000111001111011001111" & 
    "11111111111111110110110011111111001" & 
    "00000000000100000010010010111110010" & 
    "00000000000111010000110010101110111" & 
    "00000000001001011000111000101100111" & 
    "00000000001001100010101011010000100" & 
    "00000000000110000011011111100010001" & 
    "11111111111111000001110100110010001" & 
    "11111111111000011010100010001010010" & 
    "11111111110110010111000000110110001" & 
    "11111111111001100011110010100100011" & 
    "11111111111011100100110011010000100" & 
    "11111111111001111000000111111011111" & 
    "11111111110111110011001111010000110" & 
    "11111111111000001010111101111010001" & 
    "11111111111110001001111110010001001" & 
    "00000000000101100110000001111111101" & 
    "00000000001010000111000010100110000" & 
    "00000000001001001101101101000010001" & 
    "00000000000011100010000000011001101" & 
    "11111111111110001100100110110010101" & 
    "11111111111011010010011011011110011" & 
    "11111111111001110011011110011011110" & 
    "11111111110110111101010000111111100" & 
    "11111111110010100011111011111100100" & 
    "11111111101111111100110101001100000" & 
    "11111111110010000100110000000101111" & 
    "11111111111011110010000010000000101" & 
    "00000000001000000001001000010111110" & 
    "00000000001111000010100101010100001" & 
    "00000000001101000001111100100111011" & 
    "00000000000100100100011110010110110" & 
    "11111111111101000101000001010001011" & 
    "11111111111011001100011001100111011" & 
    "11111111111011100001111100011000001" & 
    "11111111111011011111100100011010011" & 
    "11111111111011110101111000000111101" & 
    "11111111111100010000101000111000000" & 
    "11111111111100110101000110101000101" & 
    "11111111111110100001101011001000011" & 
    "00000000000010001100110110100000101" & 
    "00000000000111011101010101011001100" & 
    "00000000001100110001111000001110101" & 
    "00000000001100111110011010000110001" & 
    "00000000000110011101001010001000011" & 
    "11111111111111110001011011100001001" & 
    "11111111111011111111111011000110001" & 
    "11111111111011010101010001111100100" & 
    "11111111111011111001010010110111001" & 
    "11111111111010111000111110010111110" & 
    "11111111111001101011000010101110110" & 
    "11111111111000110111111111101110011" & 
    "11111111111010001111100000111000011" & 
    "11111111111111010010001111000100111" & 
    "00000000000110010111100010010100001" & 
    "00000000001011100110011110110000011" & 
    "00000000001100011000110110100000010" & 
    "00000000001001001111011110110101000" & 
    "00000000000011100000101010111101001" & 
    "11111111111100100000000100101000000" & 
    "11111111110110011110110111100000111" & 
    "11111111110011000001111111000001110" & 
    "11111111110010110101110110000000011" & 
    "11111111110100011011101001011101011" & 
    "11111111110111111111110000100100010" & 
    "11111111111110001111110000100001100" & 
    "00000000000011101101000010100011110" & 
    "00000000000110101011001011110101011" & 
    "00000000000110111101101111011001110" & 
    "00000000000011000001001111001000011" & 
    "11111111111110100111110011011110010" & 
    "11111111111110110011101111001101011" & 
    "00000000000010100001101000100100110" & 
    "00000000000101010011001000000001011" & 
    "00000000000001011010001001010011011" & 
    "11111111111001101110001001011011101" & 
    "11111111110111010110101110101111000" & 
    "11111111111111000000111111000100011" & 
    "00000000001001110010010001110011101" & 
    "00000000001110110111011000001000001" & 
    "00000000001101010101100111100000111" & 
    "00000000001000000011100010100100110" & 
    "00000000000011011010010111001000001" & 
    "00000000000000001110110100001011100" & 
    "11111111111010111010011001001100101" & 
    "11111111110101100100110010001111001" & 
    "11111111110001100100001110100110010" & 
    "11111111110000000110111110100011100" & 
    "11111111110010000001111100011110011" & 
    "11111111110111001011111100101011001" & 
    "11111111111111000100101000110100100" & 
    "00000000000111100100010011110000001" & 
    "00000000001101010011100100010000110" & 
    "00000000001100111010011000000100001" & 
    "00000000000110000001011010000000100" & 
    "11111111111101001111011101100110100" & 
    "11111111110111100111110011110111001" & 
    "11111111110111011111000010001011011" & 
    "11111111111010001100100110000001101" & 
    "11111111111011101100100110111001111" & 
    "11111111111101001011011111000100000" & 
    "00000000000000111001101101000110101" & 
    "00000000000110001001011001001101101" & 
    "00000000001001000111011100111011001" & 
    "00000000000110010000011101001100000" & 
    "00000000000010010010101111010111000" & 
    "00000000000010000100011001010111100" & 
    "00000000000100011100111101000000101" & 
    "00000000000101001010010100011000000" & 
    "11111111111111111110101011000100010" & 
    "11111111110111111111111110101000101" & 
    "11111111110010000010011011101011000" & 
    "11111111110001000100100011010000010" & 
    "11111111110100011001011100110010100" & 
    "11111111111001111001111100110111101" & 
    "00000000000000001000101010100001001" & 
    "00000000000101100010111011100010000" & 
    "00000000001010000000101011010110010" & 
    "00000000001110011101101011010110001" & 
    "00000000010000001111010100011101001" & 
    "00000000001101101111001100110101000" & 
    "00000000000110100011111110110010101" & 
    "11111111111101101111111011001010010" & 
    "11111111111001011011011111110001101" & 
    "11111111111001110111000011000011001" & 
    "11111111111011000110100010011011010" & 
    "11111111111000100001010010001100000" & 
    "11111111110011100101111100101010111" & 
    "11111111110100110101000101000111001" & 
    "11111111111101110011110101001010100" & 
    "00000000001001010001010010100110000" & 
    "00000000001111001001111010000000100" & 
    "00000000001101001000011001000000101" & 
    "00000000000110110010100000111011100" & 
    "11111111111110010101010011110011011" & 
    "11111111110111111011111110001001101" & 
    "11111111110101000000011111100101110" & 
    "11111111110111011010100100101111110" & 
    "11111111111101111001110000100110000" & 
    "00000000000011001001001100101110100" & 
    "00000000000111011001010111000011111" & 
    "00000000001001101100000101000001111" & 
    "00000000000111110000001101100000010" & 
    "00000000000010111000101011110100101" & 
    "11111111111110101011011111100010010" & 
    "11111111111110100010100010010001100" & 
    "11111111111110011110101010010110011" & 
    "11111111111011011111011111110100110" & 
    "11111111110101110001000010011011001" & 
    "11111111110010010000110001100001110" & 
    "11111111110100001011011011001000000" & 
    "11111111111001100011001110100101111" & 
    "00000000000000001011000001010110100" & 
    "00000000000110111110100110010111110" & 
    "00000000001010100001101111001110111" & 
    "00000000001000111111110101100001100" & 
    "00000000000011011001000001011110000" & 
    "11111111111101010011101000001011001" & 
    "11111111111010100100100000001011110" & 
    "11111111111011011111101110100111111" & 
    "11111111111101010000101011101000111" & 
    "11111111111100101110000000101010010" & 
    "11111111111010100101111010001001010" & 
    "11111111111011001111010011111101110" & 
    "11111111111111000001111001010001110" & 
    "00000000000101010011011000100110010" & 
    "00000000001001011101011000000101001" & 
    "00000000001010000111010110100011011" & 
    "00000000001001011001111011101101101" & 
    "00000000000110110010010010100011001" & 
    "00000000000010101110011000100101110" & 
    "11111111111110000000110111001011001" & 
    "11111111111001011110110001111100011" & 
    "11111111110110001110010101110011010" & 
    "11111111110101111011111011100010010" & 
    "11111111111001100100111100110110100" & 
    "11111111111110100111110111100101110" & 
    "00000000000011000111110001100011111" & 
    "00000000000101100011001001011011100" & 
    "00000000000110100111110110100111111" & 
    "00000000001000011010100100111000110" & 
    "00000000001000101110101100110111110" & 
    "00000000000110001111011100111001001" & 
    "00000000000010000011001001000001101" & 
    "11111111111110101010010101110010100" & 
    "11111111111110011011100101110010001" & 
    "11111111111111010011010011111101100" & 
    "11111111111100101110000100110000000" & 
    "11111111110111001011100110100001100" & 
    "11111111110100100001101000110011011" & 
    "11111111111001101101000110001011111" & 
    "00000000000100001000100100111010111" & 
    "00000000001100011111011010111000111" & 
    "00000000001110100011000101010111100" & 
    "00000000001011010111011000101001010" & 
    "00000000000110111110100101111010101" & 
    "00000000000001011001101111100001101" & 
    "11111111111100111000001111110010010" & 
    "11111111111101110110110000000011111" & 
    "00000000000000011101110110000001110" & 
    "11111111111111001010101011000110011" & 
    "11111111111000110100110110111100000" & 
    "11111111110011010001001101101010101" & 
    "11111111110101001100101101111000101" & 
    "11111111111100110111011110100100000" & 
    "00000000000100001100100110010111101" & 
    "00000000000110110101101111011111000" & 
    "00000000000110010000111011100101100" & 
    "00000000000100011110100110101100111" & 
    "00000000000011110000110100011011111" & 
    "00000000000101011010101011000100111" & 
    "00000000000011010010001001111011001" & 
    "11111111111011101100111110001010101" & 
    "11111111110011111011101101100101010" & 
    "11111111110001100001111000000100000" & 
    "11111111110110001110100111000011101" & 
    "11111111111110011011010011101001001" & 
    "00000000000111001100100111110011110" & 
    "00000000001110001000110111011010100" & 
    "00000000001111001111001100101001110" & 
    "00000000001001010111111110000100100" & 
    "00000000000000110000010000001011101" & 
    "11111111111011111100010001100000001" & 
    "11111111111001110011100010101011100" & 
    "11111111110110111010111001101100111" & 
    "11111111110100110000110011110110011" & 
    "11111111110100101111101100010000100" & 
    "11111111110111011001110100100111110" & 
    "11111111111101001000001011000101101" & 
    "00000000000011010001101111110110100" & 
    "00000000001000011111001110000011100" & 
    "00000000001010001101100111110101001" & 
    "00000000001000001100010010100111001" & 
    "00000000000100100000000001100010110" & 
    "00000000000000100010000001100100111" & 
    "11111111111101011111010110111011111" & 
    "11111111111100000100011110111100001" & 
    "11111111111100110000000101010101010" & 
    "11111111111100110111101101101011011" & 
    "11111111111011000010001110001100101" & 
    "11111111111010101100010101011000111" & 
    "11111111111100111010110000100101010" & 
    "00000000000001100101011011110010010" & 
    "00000000000101110100011100110111011" & 
    "00000000000111101001100000011101001" & 
    "00000000000111001011011101010000001" & 
    "00000000000100010011100010001010010" & 
    "11111111111111110111000000100001100" & 
    "11111111111011001000010111111001101" & 
    "11111111111000001001111000010010100" & 
    "11111111111001001011100000001011100" & 
    "11111111111011110000110101010000010" & 
    "11111111111110100001000100001100001" & 
    "00000000000011010101101001000001011" & 
    "00000000001001101111001100110100010" & 
    "00000000001111001000010101110000110" & 
    "00000000001111010110010001101010101" & 
    "00000000001000111011100100001110001" & 
    "00000000000010101111100100000110001" & 
    "11111111111111111111110110010110111" & 
    "11111111111101100111101101101011001" & 
    "11111111111001111001110101011100111" & 
    "11111111111000001100100000010111100" & 
    "11111111111011101011101001101001001" & 
    "00000000000011001111000001011111010" & 
    "00000000001011010101101100001111110" & 
    "00000000001100110011101111101111101" & 
    "00000000000110101000100100111101101" & 
    "11111111111110111111000100001000010" & 
    "11111111111011000101101010111111011" & 
    "11111111111110100000011110010101011" & 
    "00000000000010111111101111110101111" & 
    "00000000000010001000011011100011100" & 
    "11111111111100111000100010111000110" & 
    "11111111110110100101100100000000001" & 
    "11111111110010101001001110001110010" & 
    "11111111110001111101011111101000101" & 
    "11111111110110101100011000111010111" & 
    "11111111111111010111000001011011001" & 
    "00000000000110001000100111110101010" & 
    "00000000001000001101101111111011111" & 
    "00000000000101001000011000100010101" & 
    "00000000000000101101101000111011000" & 
    "11111111111110000111110100010110100" & 
    "11111111111100100101001101000011100" & 
    "11111111111011111000001010101101001" & 
    "11111111111011101101100100000001001" & 
    "11111111111011110100101100011101101" & 
    "11111111111100110010000101010011101" & 
    "11111111111111100110100110001000010" & 
    "00000000000100011111001100010000010" & 
    "00000000001001111111001100111110000" & 
    "00000000001110111000101001110001010" & 
    "00000000001111111100111000110001111" & 
    "00000000001100101001101000001001110" & 
    "00000000001000100011011100100100100" & 
    "00000000000011111011100111111101000" & 
    "11111111111111000000100010011011101" & 
    "11111111111010101100111100010011100" & 
    "11111111111000000100100100110000101" & 
    "11111111111010001111010111110111100" & 
    "00000000000001000011111000111111101" & 
    "00000000000111001000000110110110110" & 
    "00000000001001110110001001001111010" & 
    "00000000001001000111111011111110001" & 
    "00000000000110001101010000011000010" & 
    "00000000000011011100110101011101111" & 
    "00000000000010010100011101101100010" & 
    "00000000000001100001101111010011110" & 
    "00000000000000010000111000100110111" & 
    "00000000000000100100101000101010001" & 
    "00000000000001100001101110011100110" & 
    "00000000000001110111011011100001111" & 
    "00000000000010101000011011111110100" & 
    "00000000000010101100100100011010011" & 
    "00000000000010010110010000111000110" & 
    "00000000000010001011010110101110000" & 
    "00000000000011001100000000000011001" & 
    "00000000000110110110110000000111010" & 
    "00000000001010001010111001011011111" & 
    "00000000001000011111100010010001000" & 
    "00000000000001101111100101011000110" & 
    "11111111111010110011100110011011110" & 
    "11111111110111010011000111000101000" & 
    "11111111110110000100000101110101111" & 
    "11111111110110100101011010111011101" & 
    "11111111111001000000110011111101000" & 
    "11111111111101001010100000101011011" & 
    "00000000000000100100000111001111011" & 
    "11111111111111011000001011111001010" & 
    "11111111111100011111011101000111110" & 
    "11111111111011000110100000010100001" & 
    "11111111111010001100100010000110011" & 
    "11111111111001001101111101001011010" & 
    "11111111110110001011011111111110000" & 
    "11111111110010010011101000010011011" & 
    "11111111110000111010011100100001010" & 
    "11111111110011011111110110111001010" & 
    "11111111111001010111011100000111000" & 
    "11111111111111110111001010011101011" & 
    "00000000000100010111001010111001100" & 
    "00000000000011111001001101010001111" & 
    "00000000000000110101101110010100100" & 
    "00000000000001111101001010010100100" & 
    "00000000000111101011100001111001111" & 
    "00000000001100001100000011011111110" & 
    "00000000000111101111000111011101010" & 
    "11111111111100001100111000110101001" & 
    "11111111110100001000101011110001111" & 
    "11111111110010110101010100001010011" & 
    "11111111110110111101111011001111111" & 
    "11111111111011111001011001101010000" & 
    "11111111111111001110011001010011000" & 
    "00000000000001011101000001011111111" & 
    "00000000000000101110101010111000001" & 
    "11111111111110110111011001010101010" & 
    "11111111111111011011001011101110010" & 
    "00000000000001111111001111001100110" & 
    "00000000000010001000110001111101000" & 
    "11111111111110001111110110011111110" & 
    "11111111111011101000010101110011000" & 
    "11111111111010110001101111110100100" & 
    "11111111111011001111001001010011011" & 
    "11111111111011101100011000001101011" & 
    "11111111111101011111010111000000111" & 
    "00000000000100100100000110110011100" & 
    "00000000001110100110111111100110010" & 
    "00000000010101111111011010001110000" & 
    "00000000010110010000111001010101111" & 
    "00000000001110100001010011010000101" & 
    "00000000000011110001000000000010111" & 
    "11111111111001111100010111000001010" & 
    "11111111110100011001010000000101011" & 
    "11111111110100000010110000010111001" & 
    "11111111110101111011100000101111001" & 
    "11111111110111011001000100001100001" & 
    "11111111110111110100100001011001011" & 
    "11111111111001111010100001011110000" & 
    "11111111111111000010100111011001110" & 
    "00000000000100100000101111010010111" & 
    "00000000000111001001100010100001000" & 
    "00000000000110110010001110011010101" & 
    "00000000000110100001101100000101101" & 
    "00000000000110110111011000010101010" & 
    "00000000000100010100110111100000001" & 
    "11111111111101000101101001111001101" & 
    "11111111110011110110111110111010011" & 
    "11111111101110110000100000011010100" & 
    "11111111110001101101001000111010100" & 
    "11111111111000110011101111010110001" & 
    "00000000000000000011001111001010100" & 
    "00000000000101100101011011111011110" & 
    "00000000001010001001100010010011011" & 
    "00000000001110011010111010010001000" & 
    "00000000001110001001010000011100001" & 
    "00000000001000100100101111110010110" & 
    "00000000000001110010100011001001001" & 
    "11111111111110001000110101011101110" & 
    "11111111111100011110001010100110101" & 
    "11111111111000010001010101011110100" & 
    "11111111110010100110101111001101100" & 
    "11111111101111001010110000011001110" & 
    "11111111110010011110110111010011011" & 
    "11111111111011100101010011111000011" & 
    "00000000000011000001101101101111001" & 
    "00000000000101011000101111001100000" & 
    "00000000000100010100110100100011110" & 
    "00000000000010110000000100001001111" & 
    "00000000000010111010001110011111011" & 
    "00000000000010000100110111100100100" & 
    "11111111111110010111100011101110010" & 
    "11111111111001010111011111000010101" & 
    "11111111110111100010111000001110111" & 
    "11111111111010001010111000110100111" & 
    "11111111111101111001010011001011000" & 
    "00000000000010000001101001101011011" & 
    "00000000000100111011100111111011001" & 
    "00000000000101000110101110101000110" & 
    "00000000000011111000100111011100010" & 
    "00000000000001110010000111011101111" & 
    "00000000000000111001101000011010011" & 
    "11111111111111100011001000000000001" & 
    "11111111111100100011011011110100110" & 
    "11111111110111011110011001010011011" & 
    "11111111110001000011110111000100000" & 
    "11111111101100110001111010110010101" & 
    "11111111101011110101111010100001100" & 
    "11111111101111011111100111101000101" & 
    "11111111110110111010100010100001111" & 
    "11111111111111000101110000001011101" & 
    "00000000000111001010111100110011010" & 
    "00000000001100110110111010010010100" & 
    "00000000001100110011100100111010011" & 
    "00000000000101011010101001101110011" & 
    "11111111111010000011111110001101111" & 
    "11111111110000111010011001111100000" & 
    "11111111101101111010100001000110110" & 
    "11111111110001110000111110100110001" & 
    "11111111111010001110011101100100100" & 
    "00000000000000011110010100110101011" & 
    "00000000000000101101001011000101110" & 
    "11111111111111101111011111011100000" & 
    "00000000000100111001010001111000100" & 
    "00000000001101111001010100111111100" & 
    "00000000010000101110111110110011000" & 
    "00000000001010111110011100001000101" & 
    "00000000000000111011111010011010001" & 
    "11111111111010011011110110110000010" & 
    "11111111111001100101000101101010011" & 
    "11111111110111111100011110100100111" & 
    "11111111110100011001000001110100101" & 
    "11111111110010101100001001001001101" & 
    "11111111110110001100001101000110001" & 
    "11111111111110100100100011101001111" & 
    "00000000000111011010100001011110111" & 
    "00000000001101001011100101101010111" & 
    "00000000001110010011100110111001000" & 
    "00000000001100001111111111001001011" & 
    "00000000000111111100010101110011001" & 
    "00000000000001111001011111011010010" & 
    "11111111111100001010001111110000010" & 
    "11111111110111000111000001000000011" & 
    "11111111110100000001110110111001000" & 
    "11111111110101011000010110001000001" & 
    "11111111111011000111000001110001100" & 
    "00000000000001000110101010111011100" & 
    "00000000000010010111110110010000001" & 
    "00000000000000100101011100000011110" & 
    "00000000000000101110000111110001111" & 
    "00000000000011011110000111001101110" & 
    "00000000000111100011011011111100111" & 
    "00000000001001010100110100100010000" & 
    "00000000000101110011011000011010000" & 
    "11111111111101100010011110110100110" & 
    "11111111110010100110101011110001011" & 
    "11111111101101101001100001001000000" & 
    "11111111110101000111100101000011011" & 
    "00000000000011101110110011100001111" & 
    "00000000001111000111101011000010011" & 
    "00000000010000110111011000010000000" & 
    "00000000001011010010000010101001100" & 
    "00000000000100001010011111100110110" & 
    "11111111111111100001000010010011011" & 
    "11111111111100010000001111111000000" & 
    "11111111111001101100000110101101001" & 
    "11111111111010000101010011101100000" & 
    "11111111111100110000110100010111011" & 
    "11111111111110111010001100001000100" & 
    "11111111111110011000100110011011110" & 
    "11111111111100001011101001110010001" & 
    "11111111111111101101010111000000101" & 
    "00000000001001001011110110000100001" & 
    "00000000001111101001001110100110001" & 
    "00000000001101000000000110110100011" & 
    "00000000000011110010001101000000111" & 
    "11111111111101011001100101100001010" & 
    "11111111111101010101100110110101001" & 
    "11111111111110101000111010101111011" & 
    "11111111111101011101000000000111110" & 
    "11111111111001001000110110111000010" & 
    "11111111110110011111000100110001101" & 
    "11111111110111101000001100101001001" & 
    "11111111111011010010100010110001110" & 
    "11111111111111011010010111110001101" & 
    "00000000000001111110101101110101101" & 
    "00000000000100001111100000010001101" & 
    "00000000000110101000101011110000100" & 
    "00000000000110111001111011000100000" & 
    "00000000000011001110001011101101000" & 
    "11111111111100111011001100100000011" & 
    "11111111111000100000100110100101001" & 
    "11111111110101110000001100111000000" & 
    "11111111110101100011100110100011011" & 
    "11111111110111010110110000010111001" & 
    "11111111111000100110111111001010101" & 
    "11111111111010111000011100010101111" & 
    "11111111111101011101100001111100110" & 
    "00000000000000010010111000011001111" & 
    "00000000000011011110100101100011110" & 
    "00000000000100010101100100010011110" & 
    "00000000000011010110110101111101000" & 
    "00000000000001100000110010100101010" & 
    "11111111111111010011011100001011110" & 
    "11111111111100110100111010100001000" & 
    "11111111111010100001101010100101011" & 
    "11111111111010110111010000011100101" & 
    "11111111111100110111111100101001100" & 
    "11111111111111110100010111011101111" & 
    "00000000000011100100001110111010101" & 
    "00000000000101010110011100100111110" & 
    "00000000000100111000111100101101101" & 
    "00000000000010110101001001110001100" & 
    "00000000000001111000101000000010000" & 
    "00000000000011000111000100011111000" & 
    "00000000000011100000011000100101100" & 
    "11111111111110011000101010000010110" & 
    "11111111110011011000101010000000110" & 
    "11111111101011101100000011100111010" & 
    "11111111101100111111101000100110010" & 
    "11111111110101110111011100011100010" & 
    "00000000000001001011101100011011000" & 
    "00000000000110000110110100001001111" & 
    "00000000000100010100110001111001010" & 
    "00000000000011101011000101100011011" & 
    "00000000000110110101001100111101111" & 
    "00000000001000001110111100101100010" & 
    "00000000000001101001111100110101000" & 
    "11111111110100101111100100101001111" & 
    "11111111101100011110100111000100000" & 
    "11111111101111111001101001100111111" & 
    "11111111111001100110111000100110101" & 
    "11111111111111110110100111010011110" & 
    "00000000000000111010011111110111110" & 
    "00000000000000110010000100110010101" & 
    "00000000000001011001001101000001101" & 
    "00000000000010001100001111000011110" & 
    "00000000000001010011000111111110111" & 
    "11111111111110110000111101001001011" & 
    "11111111111100001111011101000011110" & 
    "11111111111001001100001001111011001" & 
    "11111111110110011110011000011010110" & 
    "11111111110100001000100000001110000" & 
    "11111111110011000000000001001011010" & 
    "11111111110110001001000101000000000" & 
    "11111111111101110011101001011000111" & 
    "00000000000110111001000000000101001" & 
    "00000000001011001010101100111100011" & 
    "00000000000101111000101011110010111" & 
    "11111111111100100011110001110010101" & 
    "11111111111001010000101100100111001" & 
    "00000000000000000010000000010101100" & 
    "00000000001000010010001100010011111" & 
    "00000000000111001000100000101100010" & 
    "11111111111011101100100010000010111" & 
    "11111111110001101110001011001101110" & 
    "11111111110011100001101110110111010" & 
    "11111111111011101111010001110110111" & 
    "00000000000001011000110000011001000" & 
    "00000000000001111100011010101100000" & 
    "11111111111111111000100011011001010" & 
    "11111111111111110101011011011010011" & 
    "00000000000010010011010101110010010" & 
    "00000000000101001101100001110100010" & 
    "00000000000111010101111001110011000" & 
    "00000000000101110000111101000101111" & 
    "11111111111111010101011110010100100" & 
    "11111111110110110001011111010010110" & 
    "11111111110000010010010100000011001" & 
    "11111111110000100111000001011110101" & 
    "11111111110111110110011110011001001" & 
    "00000000000010000100000000111011110" & 
    "00000000001001010111001111110100110" & 
    "00000000001010000010110111010100000" & 
    "00000000000111110000100010011010011" & 
    "00000000000110110010111101010010000" & 
    "00000000000111110011010101111101111" & 
    "00000000000100111110101100011000010" & 
    "11111111111100111100100111111000010" & 
    "11111111110100111111001110000010100" & 
    "11111111110001000110010111001001000" & 
    "11111111110010100100100111011000010" & 
    "11111111110110111001000100100101100" & 
    "11111111111101000111110001101010110" & 
    "00000000000101101101010110011111010" & 
    "00000000001011101001110111011010100" & 
    "00000000001010101111001111111111001" & 
    "00000000000011001100011111101011100" & 
    "11111111111010100000100001001010010" & 
    "11111111110101100011110001101111001" & 
    "11111111110100010010000011111101110" & 
    "11111111110111111000001010001001110" & 
    "11111111111110011111101101100011011" & 
    "00000000000011000011111000100000001" & 
    "00000000000011000000010000111010000" & 
    "11111111111111111101010011111100000" & 
    "00000000000000011101101100000011010" & 
    "00000000000110100111101100110110010" & 
    "00000000001101001110100010111010101" & 
    "00000000001110000011111001100100100" & 
    "00000000001000111100110010111111000" & 
    "00000000000011010011000100110011111" & 
    "11111111111101101111100011001110011" & 
    "11111111111000111110101010011000010" & 
    "11111111110111001100000111010010101" & 
    "11111111110110110001011011000010111" & 
    "11111111110110011100001111010010010" & 
    "11111111110110111000110100010110001" & 
    "11111111111010111110110011000100101" & 
    "00000000000100101110110101010001000" & 
    "00000000001100111011110110110011000" & 
    "00000000001101110100000010101111001" & 
    "00000000001001010001100010000010001" & 
    "00000000000110101101010110010000000" & 
    "00000000000110010000100111011101110" & 
    "00000000000010001111010100011011100" & 
    "11111111111100011001010001101000010" & 
    "11111111111000100001110100010100001" & 
    "11111111110111111011100110110000110" & 
    "11111111111001000101100011101110101" & 
    "11111111111001111100111110011010110" & 
    "11111111111101001010000111101101011" & 
    "00000000000010101010111011001001110" & 
    "00000000000111010101100001000010011" & 
    "00000000000111001101011000100111000" & 
    "00000000000010100011101110101111011" & 
    "11111111111111101100111011101011011" & 
    "11111111111111011010111001000100110" & 
    "11111111111111010010011001111111101" & 
    "11111111111110111101011010100100001" & 
    "11111111111111011101001000101100011" & 
    "00000000000010010000101111010001000" & 
    "00000000000011111001111000010110110" & 
    "00000000000010100010001011001010000" & 
    "00000000000001011000111010101010100" & 
    "00000000000010101111010001110010000" & 
    "00000000000101111000010110001000100" & 
    "00000000000110011101010110000011111" & 
    "00000000000101100011000001000111001" & 
    "00000000000101100000010101110011110" & 
    "00000000000100101110011001100000110" & 
    "00000000000000101111011011100011110" & 
    "11111111111010011001110100101110010" & 
    "11111111110110000111101011001110100" & 
    "11111111110110011100111101111101111" & 
    "11111111111011001010101100100010110" & 
    "00000000000011001001101100110010101" & 
    "00000000001001111010101100010000100" & 
    "00000000001011011001100111111000110" & 
    "00000000001010011100110011110011111" & 
    "00000000001011101110100101110010110" & 
    "00000000001101110010010101011101010" & 
    "00000000001010011110001111001000001" & 
    "00000000000001101110001011100101110" & 
    "11111111111001011111111001100110111" & 
    "11111111110111000001101100100101100" & 
    "11111111111011110110110110110101110" & 
    "00000000000010110000100110110101001" & 
    "00000000000111111101110000000101100" & 
    "00000000001011010000111111110011000" & 
    "00000000001000110111101110000101011" & 
    "00000000000010100100001001000110001" & 
    "11111111111101010000111111100111101" & 
    "11111111111010110011110000001100110" & 
    "11111111111001111010100111100001101" & 
    "11111111111001010111100110111001001" & 
    "11111111111010101010101100001001000" & 
    "11111111111110001100010010001011011" & 
    "00000000000001010010110101001011001" & 
    "00000000000010100111001101011110101" & 
    "00000000000001101101111101001100111" & 
    "00000000000001111110110111101001111" & 
    "00000000000100011010010110011111010" & 
    "00000000000111010010100100000000000" & 
    "00000000000111001110010000000110101" & 
    "00000000000100010001010100100110011" & 
    "00000000000001110010011110000001100" & 
    "11111111111110011011001010111100000" & 
    "11111111111001110100011110110101000" & 
    "11111111110101110110011011101001011" & 
    "11111111110011110001100100001100110" & 
    "11111111110110000100110011000101111" & 
    "11111111111011110001000010100010000" & 
    "00000000000000011011010100000100101" & 
    "00000000000000100010010111110000011" & 
    "11111111111110110011101101010100011" & 
    "00000000000001001001001001100010000" & 
    "00000000001000100001111100100000010" & 
    "00000000001111011001111110111001100" & 
    "00000000001110011111000000011101100" & 
    "00000000000101001000011111110010000" & 
    "11111111111100000100100001111001010" & 
    "11111111111000011010011011000000011" & 
    "11111111110111100101101011111101001" & 
    "11111111111000000000000001111010110" & 
    "11111111111000101110110001100000010" & 
    "11111111111010110101001101111011101" & 
    "00000000000000110111100000011000000" & 
    "00000000001001110101101111000111100" & 
    "00000000010000111110100110001000000" & 
    "00000000001111010101011001100001001" & 
    "00000000000101010011101111000101001" & 
    "11111111111011110110001001101011100" & 
    "11111111111001000111100000101111101" & 
    "11111111111011101011001110111111100" & 
    "11111111111100101001011000000011010" & 
    "11111111111010111010001001101010001" & 
    "11111111111010011010111111110100100" & 
    "11111111111101000101101110011110001" & 
    "00000000000010011111011111001110010" & 
    "00000000001001010100110010000110110" & 
    "00000000010011011001101011100110001" & 
    "00000000011001101100111100101111010" & 
    "00000000010100011110101110100000111" & 
    "00000000000110101001010110000010101" & 
    "11111111110111101110111001000110010" & 
    "11111111110000001000111100101110011" & 
    "11111111101110011100000101001010110" & 
    "11111111101111110111010110101011111" & 
    "11111111110101111001000001110111101" & 
    "11111111111110011101100101000000010" & 
    "00000000000101000011011001011101101" & 
    "00000000000111011011101101011101111" & 
    "00000000001001000110001110101001011" & 
    "00000000001100100011010110001011101" & 
    "00000000001111001110011101010000111" & 
    "00000000001101011100101101001011000" & 
    "00000000000111001001101101111101001" & 
    "00000000000000101000010010101100111" & 
    "11111111111010110111011001111111011" & 
    "11111111110101111000110001011001100" & 
    "11111111110101000010010111011101110" & 
    "11111111111000011001001011000101011" & 
    "11111111111101011101000110010111010" & 
    "00000000000010111111100001011101010" & 
    "00000000000111101010100000110000000" & 
    "00000000001011010110111010010110000" & 
    "00000000001100111011101011000100100" & 
    "00000000001011001001011100101111000" & 
    "00000000000101101011110000010111011" & 
    "11111111111101110100110000001010100" & 
    "11111111111000101110101111100001100" & 
    "11111111110111100010001110000110110" & 
    "11111111111010000000010100110011111" & 
    "11111111111111010001001101010010111" & 
    "00000000000011111100111011100001101" & 
    "00000000000110110011111011010111000" & 
    "00000000000111000111010000110000010" & 
    "00000000000100101110100110010010011" & 
    "00000000000000101000000100001001000" & 
    "11111111111110010011011010111001101" & 
    "00000000000000001101100100010010101" & 
    "00000000000010110001011101000110010" & 
    "00000000000100111111001001111000000" & 
    "00000000000100011011010001101110011" & 
    "11111111111110100011100111010101111" & 
    "11111111110111000110100100100101011" & 
    "11111111110100101000110010111100000" & 
    "11111111111010000010011100111100011" & 
    "00000000000010010110100001100000001" & 
    "00000000000110001011010101010111000" & 
    "00000000000100110101111011000100011" & 
    "00000000000011111011100110011111101" & 
    "00000000000110011100010000011111100" & 
    "00000000000101110000111001100111001" & 
    "11111111111101010010010000001000101" & 
    "11111111110011011101000100110101011" & 
    "11111111110010010010000010010001000" & 
    "11111111111010011111010011000101000" & 
    "00000000000011001101111110011011010" & 
    "00000000000011000001110111100100010" & 
    "11111111111100011100111100010111010" & 
    "11111111111000010000111111110000001" & 
    "11111111111100001011010100111010000" & 
    "00000000000101010011000110110010010" & 
    "00000000001001010111101011001111110" & 
    "00000000000011111011011101010001011" & 
    "11111111111010100111010100000100101" & 
    "11111111110101111111110110010011110" & 
    "11111111110111100101001101001110011" & 
    "11111111111001011110111011011001101" & 
    "11111111110111110100111000001100110" & 
    "11111111110011111001001110001000001" & 
    "11111111110100110011001111001101000" & 
    "11111111111101010001110101000010000" & 
    "00000000000110110100111100110111100" & 
    "00000000001010111111001001000101111" & 
    "00000000000110101000100101110010010" & 
    "11111111111110010110011001001110010" & 
    "11111111111011100010010111000111000" & 
    "11111111111110110101010100011110001" & 
    "00000000000010101010111111100100110" & 
    "00000000000001111110111100000001011" & 
    "11111111111101000100101110001101010" & 
    "11111111111000101101111101011111101" & 
    "11111111111001001010110000111000010" & 
    "00000000000000110001011100100000100" & 
    "00000000001011010101100010101110110" & 
    "00000000010010000011000010010000011" & 
    "00000000010001001001110000011001001" & 
    "00000000001010001111111110111101110" & 
    "00000000000011100111011001010001000" & 
    "11111111111110011100000101100111100" & 
    "11111111111011010111001110011010010" & 
    "11111111111010111001110011011110000" & 
    "11111111111010111100001001011011000" & 
    "11111111111100010100000101001100001" & 
    "11111111111110100001101111111000111" & 
    "00000000000000010010011010111100111" & 
    "00000000000010110110010010011011110" & 
    "00000000000110011110110010101111011" & 
    "00000000001010111001110110011100100" & 
    "00000000001100111011100110111100011" & 
    "00000000001010010000000101000100110" & 
    "00000000000011111010100000011000110" & 
    "11111111111101110001010011111000111" & 
    "11111111111010100111010111011100011" & 
    "11111111111000000001111001010011000" & 
    "11111111110110111000001001111101110" & 
    "11111111111001110100100011010000100" & 
    "00000000000001000010010001101010111" & 
    "00000000001001101100000011001110101" & 
    "00000000001101000000000001000111111" & 
    "00000000001001101010100000000101101" & 
    "00000000000101001000100000010011101" & 
    "00000000000001100101001111110001011" & 
    "11111111111110101010010010110101011" & 
    "11111111111011010000100111101100000" & 
    "11111111111000100111001111010101100" & 
    "11111111111001100001011000011111001" & 
    "11111111111100011000010100010111011" & 
    "11111111111100110111000000000111111" & 
    "11111111111011000101001000110010001" & 
    "11111111111010110010110001100110011" & 
    "11111111111100110100000111101110100" & 
    "00000000000001000000111001110000011" & 
    "00000000000111111100110000100110111" & 
    "00000000001110000100010010111101111" & 
    "00000000001110001110010110110101000" & 
    "00000000001000001110101000100101111" & 
    "11111111111111011000010111111110101" & 
    "11111111111001101010011001110100000" & 
    "11111111110111100011010100100101100" & 
    "11111111110110011101111001010011000" & 
    "11111111110111010011101000101101110" & 
    "11111111111001110000000111101010101" & 
    "11111111111111011001100101001001001" & 
    "00000000000111110011000111110001010" & 
    "00000000001101101010100110110100000" & 
    "00000000001111111101100010000110000" & 
    "00000000001110000101111010010101000" & 
    "00000000001010101010110000111110110" & 
    "00000000000101001101000000001001011" & 
    "11111111111101111111100000110001000" & 
    "11111111110111011000100010011101010" & 
    "11111111110101001111011110110100010" & 
    "11111111111001111100100001111001001" & 
    "11111111111110011100011110000110100" & 
    "00000000000001110110101001100001100" & 
    "00000000000110111100011111011101000" & 
    "00000000001001010000010100000001100" & 
    "00000000000110111000010111110110010" & 
    "00000000000000111101011001111110110" & 
    "11111111111101010001100000100011111" & 
    "11111111111101011110101100101111001" & 
    "11111111111100001000110001001111000" & 
    "11111111110110100010001110001101001" & 
    "11111111110000101010011001000010110" & 
    "11111111101111111110010010100101001" & 
    "11111111110011100111000111000100010" & 
    "11111111110110111100110100011010100" & 
    "11111111111010111000011110101000101" & 
    "11111111111111100010001010001101000" & 
    "00000000000101001010111000100010110" & 
    "00000000001011000001111011010101100" & 
    "00000000001100111100000101100001100" & 
    "00000000001000001100000100000110110" & 
    "11111111111101111000101100011011111" & 
    "11111111110101100111010000001001100" & 
    "11111111110101001101110011010100111" & 
    "11111111111001111011000101011110100" & 
    "11111111111111011101100111001010111" & 
    "00000000000001011010000010000000001" & 
    "00000000000001111000001010100110111" & 
    "00000000000010000101100000001000100" & 
    "11111111111111110010001100101110100" & 
    "11111111111101001111110000001101000" & 
    "11111111111101010101110010001001000" & 
    "00000000000001101100110100100101001" & 
    "00000000001000110001001111111101010" & 
    "00000000001010100001001110110111110" & 
    "00000000000011011000100111000110100" & 
    "11111111111001010011101001101011011" & 
    "11111111110101111000010100010101111" & 
    "11111111111010010110110110100100011" & 
    "00000000000000100100000100000011000" & 
    "00000000000100010100010000101110110" & 
    "00000000000110010101001100010101001" & 
    "00000000001010001111100011111000001" & 
    "00000000001101100000011010111010111" & 
    "00000000001011010100110101001011101" & 
    "00000000000101011010110010011111100" & 
    "11111111111110111000010101011010010" & 
    "11111111111010010100000111101001001" & 
    "11111111111001110110110111110010101" & 
    "11111111111011110011000101110110101" & 
    "11111111111101000000110100111001010" & 
    "11111111111011100110101010111001010" & 
    "11111111111001011110011110100000101" & 
    "11111111111011010111100111010110110" & 
    "00000000000001110000111001110111011" & 
    "00000000001010011111111100101110010" & 
    "00000000001111111010110111000110001" & 
    "00000000001100101001101110110100101" & 
    "00000000000010111001101111110100111" & 
    "11111111110111110000110001010010111" & 
    "11111111110010000000001000011100111" & 
    "11111111110100001111000100010111010" & 
    "11111111111010101010101011011111001" & 
    "11111111111111111000000111010011111" & 
    "00000000000010001011001100010001110" & 
    "00000000000100101100111010011010101" & 
    "00000000001000011100110010111110100" & 
    "00000000001101100111001010100001001" & 
    "00000000010001100010101101011001101" & 
    "00000000010000011000110101111011111" & 
    "00000000001100010001110111000000010" & 
    "00000000000110010110001010110100101" & 
    "11111111111111001110111110000101101" & 
    "11111111111010000001110010001010010" & 
    "11111111110110101001011100111110110" & 
    "11111111110110011010111000000010110" & 
    "11111111111001100010110101101111111" & 
    "00000000000000011100000110100101010" & 
    "00000000001001110111100010110000000" & 
    "00000000010000011100101111101101110" & 
    "00000000010000110101101000100001011" & 
    "00000000001101101101111000010100111" & 
    "00000000001101011110101010101110011" & 
    "00000000001110101010010010111111000" & 
    "00000000001011001110111010010101000" & 
    "00000000000010010110100111000101110" & 
    "11111111110111101000101110000010100" & 
    "11111111110001110000011011110001001" & 
    "11111111110010101101111111000111000" & 
    "11111111111001011100101100001001010" & 
    "00000000000100000001101111000101000" & 
    "00000000001101110100100100011001100" & 
    "00000000010001010001100111011001001" & 
    "00000000001101110001100100010000000" & 
    "00000000001000101000000010010111111" & 
    "00000000000110111110000100011011001" & 
    "00000000000111001000011100110010101" & 
    "00000000000011111010110010011001001" & 
    "11111111111100100000001011011000101" & 
    "11111111110100111001100000001000111" & 
    "11111111110101010110111101101001101" & 
    "11111111111110111111111101111011001" & 
    "00000000001001111011001011011101010" & 
    "00000000001110000011111101011100000" & 
    "00000000001011001101110111101001010" & 
    "00000000001000101001010011000010010" & 
    "00000000001000000000011110100100011" & 
    "00000000000111001001000010010010101" & 
    "00000000000101001101110111100000011" & 
    "00000000000011011111100000100000010" & 
    "00000000000010111010011010011101010" & 
    "11111111111111111110111110010100110" & 
    "11111111111011001111000011111011000" & 
    "11111111111000111000101011000111100" & 
    "11111111111011001100011110000111100" & 
    "11111111111111010010110000000110010" & 
    "00000000000010000100010111110000101" & 
    "00000000000011111000010101100101100" & 
    "00000000000100111111001010011011011" & 
    "00000000000101101111010010000101111" & 
    "00000000000110101110110010110100001" & 
    "00000000000110011101111100001101000" & 
    "00000000000010110000100010101111010" & 
    "11111111111100110000000011110001000" & 
    "11111111111000101110110101011100010" & 
    "11111111111011001101111101001101001" & 
    "00000000000001001100111110000001000" & 
    "00000000000100000011000011011111010" & 
    "00000000000011010101000100011001110" & 
    "00000000000011010100011111111100000" & 
    "00000000001000010111000000111101100" & 
    "00000000001110001010101101101111000" & 
    "00000000001101111110110100001010001" & 
    "00000000000110111110000111001111111" & 
    "11111111111101011101101101001010010" & 
    "11111111111000001110101100100001000" & 
    "11111111110110111111111110001110001" & 
    "11111111110110100011011100010001001" & 
    "11111111110110010011101010000111011" & 
    "11111111110111011000110011111000001" & 
    "11111111111011000110110111110111100" & 
    "00000000000000000110000000000001010" & 
    "00000000000101010100100111111010111" & 
    "00000000001000110001100110001101010" & 
    "00000000000111111011101111011010010" & 
    "00000000000011110001001101111000001" & 
    "11111111111110111110100100001001000" & 
    "11111111111101010001101011000001100" & 
    "11111111111110001010101000011001111" & 
    "11111111111110001101000010001111101" & 
    "11111111111110001001010111000010101" & 
    "11111111111110111100011010001001101" & 
    "11111111111111100111010010001100100" & 
    "11111111111101110011101100110100100" & 
    "11111111111001011011100101111001011" & 
    "11111111110111111011110011101100101" & 
    "11111111111011001010011111000110100" & 
    "11111111111111011100011100110001100" & 
    "00000000000000010010011100001111001" & 
    "11111111111100000111110010001111001" & 
    "11111111110110110010111110001101100" & 
    "11111111110011001100010011100100011" & 
    "11111111110100100111110001100011001" & 
    "11111111111100101001000010110010100" & 
    "00000000000110110110000111010010010" & 
    "00000000001101000011101101010110001" & 
    "00000000001011111110110001101010010" & 
    "00000000001000010000001111110110111" & 
    "00000000000101111001111111011101111" & 
    "00000000000010111010010010110100010" & 
    "11111111111110110110011001001010100" & 
    "11111111111010100011111001100111010" & 
    "11111111111000001011111100001100110" & 
    "11111111111000000001101011010101011" & 
    "11111111111000111101110110001110001" & 
    "11111111111101001011111001011110111" & 
    "00000000000011001100111010000110111" & 
    "00000000000101010110101111110111011" & 
    "00000000000001111110010011100111010" & 
    "11111111111110111110011100111010011" & 
    "00000000000010011100010011011101100" & 
    "00000000001000000111011101110110011" & 
    "00000000001001111111000100110101010" & 
    "00000000000111100000010111110101111" & 
    "00000000000011000111111000110001110" & 
    "11111111111111000001100100000010110" & 
    "11111111111001001010010101100000101" & 
    "11111111110100001101000011011101000" & 
    "11111111110101010101100001001000101" & 
    "11111111111100000111101100001001100" & 
    "00000000000100110011110111110100100" & 
    "00000000001010001110000010110000011" & 
    "00000000001011000100101110100001001" & 
    "00000000001001111101101000001011100" & 
    "00000000000111010001101000100101100" & 
    "00000000000010110010101111111000111" & 
    "11111111111101000101000000001011011" & 
    "11111111111000011111111010010000001" & 
    "11111111110111100100010100110001010" & 
    "11111111111010011111010101111110101" & 
    "11111111111111010010001001100011101" & 
    "00000000000010000001110111001010100" & 
    "00000000000010010100111011111111011" & 
    "00000000000010001101100001101100100" & 
    "00000000000011001000110110110100100" & 
    "00000000000110110001010111010011001" & 
    "00000000001001000110010110011110000" & 
    "00000000000111100010110101000010011" & 
    "00000000000101001000101011010001110" & 
    "00000000000100001101001100001110010" & 
    "00000000000100011011011001111111010" & 
    "00000000000001011100010000100000010" & 
    "11111111111010111000100011010000000" & 
    "11111111110111001100111010000010000" & 
    "11111111111001101101110111011000100" & 
    "11111111111110000101100110000101100" & 
    "11111111111111101000110010101111110" & 
    "11111111111110110101101100001001101" & 
    "00000000000001011001000000110100110" & 
    "00000000000110101111011001011110010" & 
    "00000000001000011100010000010010111" & 
    "00000000000011000111111000110101111" & 
    "11111111111010110001010110011011110" & 
    "11111111110110000010011001011000000" & 
    "11111111110100110011011100001101100" & 
    "11111111110110001000110011101100010" & 
    "11111111111001111101011000110010110" & 
    "00000000000000001100001001101010011" & 
    "00000000000101010100111011111100111" & 
    "00000000000010100001010011000101010" & 
    "11111111111100110011000000111110000" & 
    "11111111111011101011101011100000001" & 
    "00000000000000100001111111111010110" & 
    "00000000000110010100111100110000110" & 
    "00000000000100100001001010111100010" & 
    "11111111111101011111101010110001000" & 
    "11111111110111111001111010111110110" & 
    "11111111110110110111100000011110010" & 
    "11111111111000110100111101110101000" & 
    "11111111111100001010000111001101011" & 
    "11111111111111100001101110101110101" & 
    "00000000000000111001110100111001110" & 
    "00000000000001110101011110001111010" & 
    "00000000000100110010111111101101111" & 
    "00000000001001101110111000111011010" & 
    "00000000001111011001110001100010100" & 
    "00000000001111100100110001100100110" & 
    "00000000000110110101100101010010010" & 
    "11111111111001011001000100011110100" & 
    "11111111101110100111001100100100011" & 
    "11111111101101111101001110010011000" & 
    "11111111110110100001011000010111100" & 
    "00000000000000010000111110111000000" & 
    "00000000000110110000100010011001001" & 
    "00000000001000100000011101101000010" & 
    "00000000001000010110001111101010101" & 
    "00000000000111110010000011010110110" & 
    "00000000000101101000101000000100110" & 
    "00000000000010100110010011111001010" & 
    "00000000000000011010011011100110011" & 
    "00000000000000001001010100111011001" & 
    "11111111111111000111100000111010001" & 
    "11111111111101001100011001110101011" & 
    "11111111111011101110011111000101010" & 
    "11111111111100100000010000100111010" & 
    "00000000000001101100000111001110011" & 
    "00000000000110100001101010000001110" & 
    "00000000000110011001101110001100110" & 
    "00000000000100111001111001000011100" & 
    "00000000000101111000011011001111000" & 
    "00000000001000011100001011001101101" & 
    "00000000000110101101101011011101010" & 
    "11111111111110100110011001100101010" & 
    "11111111110101001101010010010110001" & 
    "11111111110000111110110100011010100" & 
    "11111111110100011000101110011010010" & 
    "11111111111010100000111111101011001" & 
    "11111111111111101010011011001101100" & 
    "00000000000011001100111111010010001" & 
    "00000000000011110110000111111101011" & 
    "00000000000010100011000111000011100" & 
    "00000000000000001110000111001100110" & 
    "11111111111101011001001001011111010" & 
    "11111111111010010110001010000000001" & 
    "11111111110111010000010100001011110" & 
    "11111111110100101111100011011101110" & 
    "11111111110010010111101110010110011" & 
    "11111111110010001100100111011111100" & 
    "11111111110101000010000101011111001" & 
    "11111111111010010011100100111100111" & 
    "00000000000000111010010110010000111" & 
    "00000000000101110100100101101011001" & 
    "00000000000110100100011101010010100" & 
    "00000000000100010101110000010101000" & 
    "00000000000000011110011110110111111" & 
    "11111111111100100110100100101111101" & 
    "11111111111001011010100011111100001" & 
    "11111111110110110100011010101101101" & 
    "11111111110011010111001010111010100" & 
    "11111111101110010100000110110110100" & 
    "11111111101011110100100010000101100" & 
    "11111111110010011010101110110100101" & 
    "00000000000001101010001110010001010" & 
    "00000000010000011000100011011001000" & 
    "00000000010011110100111110001011001" & 
    "00000000001101110010110111001011111" & 
    "00000000000111000010001010011010010" & 
    "00000000000010110111000010001011010" & 
    "11111111111110011100100111101001001" & 
    "11111111111000001011001011010101011" & 
    "11111111110001011011010010001010111" & 
    "11111111101101011100110111111101101" & 
    "11111111101111001000111111010010110" & 
    "11111111110110000111011010010110111" & 
    "11111111111111100011011000001110011" & 
    "00000000000111110101111011111001100" & 
    "00000000001001111111011100001010001" & 
    "00000000000111100001110010111101000" & 
    "00000000000110010111101110011110001" & 
    "00000000000110101001000010011011101" & 
    "00000000000101110111001101110100001" & 
    "00000000000010110110111000111111000" & 
    "11111111111101101101010111110111101" & 
    "11111111111000110001001000101000101" & 
    "11111111110100101001110001111000101" & 
    "11111111110100000011000100001110001" & 
    "11111111111001100001010111110001011" & 
    "00000000000010001110011101101010001" & 
    "00000000001000001010000110000111101" & 
    "00000000001000001010100011011110101" & 
    "00000000000111011000011100100111001" & 
    "00000000001010001111101101100101000" & 
    "00000000001100101110100101001111000" & 
    "00000000001001011001001101110001011" & 
    "00000000000000011000001010101010100" & 
    "11111111111010000000011110110111111" & 
    "11111111111001000011001011111001111" & 
    "11111111111001101100001100010011010" & 
    "11111111111010010011101111100111110" & 
    "11111111111100010010000111100100000" & 
    "00000000000001110011100000111100110" & 
    "00000000000110111110111011010001101" & 
    "00000000000111011111001101001110111" & 
    "00000000000100001101001000101110110" & 
    "00000000000001000111100100000110101" & 
    "00000000000000111000010001010110011" & 
    "11111111111111010111111000111110100" & 
    "11111111111011010100010010110101001" & 
    "11111111110111011001011010000000111" & 
    "11111111110100101111110110000010101" & 
    "11111111110010111011110111010110001" & 
    "11111111110010011011010000101011011" & 
    "11111111111001001011010010111000000" & 
    "00000000001001011100101111011110100" & 
    "00000000011010110101110011111111110" & 
    "00000000100001101000100100111011001" & 
    "00000000011001000001111110011000010" & 
    "00000000001000001010110110111000010" & 
    "11111111111010111111000010001000111" & 
    "11111111110101110011000110001001011" & 
    "11111111110110111110001001111000111" & 
    "11111111111010010100010011011100100" & 
    "11111111111011100100100110110101110" & 
    "11111111111001110010001111010100001" & 
    "11111111111000011001001001011110100" & 
    "11111111111100011000011001011100101" & 
    "00000000000100100011110101100100111" & 
    "00000000001011100001100011010110001" & 
    "00000000001110110110111011101100110" & 
    "00000000001101000011111010111111000" & 
    "00000000000111100111100101111001001" & 
    "00000000000000101101101111110111000" & 
    "11111111111001110110010011100010011" & 
    "11111111110011110111100101011100110" & 
    "11111111101110100011001010011001100" & 
    "11111111101100111010001101111101001" & 
    "11111111110001001001000101001100001" & 
    "11111111111011001110110111000001110" & 
    "00000000000110100110001111101010100" & 
    "00000000001010011010001100000101100" & 
    "00000000000110111010111010111101000" & 
    "00000000000000010001000000110011010" & 
    "11111111111010110000000111111000110" & 
    "11111111111010101000011110111000010" & 
    "11111111111110000100010110101010001" & 
    "00000000000000111001110100010100011" & 
    "00000000000000111111110101101110011" & 
    "11111111111111110111011110010000000" & 
    "11111111111110011011111010001101010" & 
    "11111111111100110001111001101010111" & 
    "11111111111101101000000001110100101" & 
    "00000000000001001101101100111011101" & 
    "00000000000111010101111010110010100" & 
    "00000000001101010101010100111100011" & 
    "00000000001101111001010111011010111" & 
    "00000000001011000001001110100010111" & 
    "00000000000101110100000011100000000" & 
    "11111111111100011110000101101111110" & 
    "11111111110010101101010101011111111" & 
    "11111111101101101111011101111010011" & 
    "11111111110000010100010111101000000" & 
    "11111111111000011111100111111111011" & 
    "00000000000010001010001000111100001" & 
    "00000000001000101001101100110001010" & 
    "00000000001000111111000000011000101" & 
    "00000000000110010010011111111101010" & 
    "00000000000011011000101110001011111" & 
    "00000000000010110111001000100010101" & 
    "00000000000010100001100001011101110" & 
    "11111111111100011101101011011111110" & 
    "11111111110011111100111111101110110" & 
    "11111111101111011110111011100111001" & 
    "11111111110001011100010101000111110" & 
    "11111111110110010010000011011111011" & 
    "11111111111010011100011110011110011" & 
    "11111111111110000001100101100101100" & 
    "00000000000000000011110011011011011" & 
    "00000000000001100111100001101000000" & 
    "00000000000011101100010010101000011" & 
    "00000000000100110001111000001101011" & 
    "00000000000100001111010111100000000" & 
    "00000000000000111000001111001011010" & 
    "11111111111011011001110000000101111" & 
    "11111111110111101101010110110010101" & 
    "11111111110110100100011110001011111" & 
    "11111111110110100011001001100100001" & 
    "11111111111000110001010011010001110" & 
    "11111111111110110010010110011000010" & 
    "00000000000111001100010101110110100" & 
    "00000000001100100010001111111100100" & 
    "00000000001100101001101100101110010" & 
    "00000000000111001001110100111011110" & 
    "00000000000000101111000110011001011" & 
    "11111111111110010110110100000001000" & 
    "11111111111110110010010010101110010" & 
    "00000000000000100110110100000010100" & 
    "11111111111111100101111100110010001" & 
    "11111111111001011000011101011100000" & 
    "11111111110001000000011011010001110" & 
    "11111111101110011001101110001011110" & 
    "11111111111000001000010111001001001" & 
    "00000000001000010010101110101111011" & 
    "00000000010011101111100011111000010" & 
    "00000000010011000011000101010110010" & 
    "00000000001010001100110000010001111" & 
    "00000000000010011101100101011111110" & 
    "11111111111111111011001100101110001" & 
    "00000000000000010101110011111101111" & 
    "11111111111111000110101111010010101" & 
    "11111111111011100001011101110011010" & 
    "11111111110111110001011110110110001" & 
    "11111111110101101100110111101100100" & 
    "11111111110111010000110101010111101" & 
    "11111111111100111101001001000001101" & 
    "00000000000011011001110001000100011" & 
    "00000000001000101111111101011000010" & 
    "00000000001100100011011001111100100" & 
    "00000000001100111110010001010011011" & 
    "00000000001001101001000010011100100" & 
    "00000000000011000111011110010010001" & 
    "11111111111100010000010011010000011" & 
    "11111111110111001010111111111000110" & 
    "11111111110011110101100101000110111" & 
    "11111111110010000000001000011010000" & 
    "11111111110011100100111000010101000" & 
    "11111111111100100011011011001110000" & 
    "00000000001001010011010101100101000" & 
    "00000000010000001010111111111101101" & 
    "00000000001101000011000111111001101" & 
    "00000000000110100010111011101100111" & 
    "00000000000110000011111110110100001" & 
    "00000000001010011111101101000100100" & 
    "00000000001001100011001001110100011" & 
    "11111111111111001011110001001010000" & 
    "11111111110011010100000001001010100" & 
    "11111111110001111111111000101010010" & 
    "11111111111010101000100101111101001" & 
    "00000000000011101010100101100110100" & 
    "00000000000110110011100000011001111" & 
    "00000000000101110101000110111001001" & 
    "00000000000110011100000000101010100" & 
    "00000000001000011100011011110100011" & 
    "00000000000111011111011010101010110" & 
    "00000000000010101110001001101110010" & 
    "11111111111101011110111101011100011" & 
    "11111111111011111010110000010001110" & 
    "11111111111011101010011000100100000" & 
    "11111111111000111111100110100011000" & 
    "11111111110100111101111101110100011" & 
    "11111111110101100110010111011101000" & 
    "11111111111101011101010110010100100" & 
    "00000000000101000000100111010101010" & 
    "00000000000100110001010001100100101" & 
    "11111111111111111010011000110101101" & 
    "11111111111110000101100001011100000" & 
    "00000000000001111100010110010011111" & 
    "00000000000010110101101101110110100" & 
    "11111111111011010011001111000101100" & 
    "11111111110010011010101010001110111" & 
    "11111111101111101001101011110100010" & 
    "11111111110100111010011100100000101" & 
    "11111111111100011001100011010101100" & 
    "00000000000001010000011010011000100" & 
    "00000000000011111001011001001010000" & 
    "00000000000110101000101001111101010" & 
    "00000000001001101110010100001000000" & 
    "00000000001001001101000111010001111" & 
    "00000000000111000101001011111111110" & 
    "00000000000101011100101111010001000" & 
    "00000000000011010101001000100110101" & 
    "00000000000000101100111110100011111" & 
    "11111111111011110001111001111111010" & 
    "11111111110110000011000011100101001" & 
    "11111111110010111101101011001110110" & 
    "11111111110101111101000010111101010" & 
    "11111111111110101011111111110010000" & 
    "00000000001000111111101010001111101" & 
    "00000000001110100101001100111111110" & 
    "00000000001100011011000100001111110" & 
    "00000000001000000101011000111101110" & 
    "00000000000110111110010000001010000" & 
    "00000000000110100111010110000011010" & 
    "00000000000010001100111110010111001" & 
    "11111111111100000110110001001001010" & 
    "11111111111001101010111111111001001" & 
    "11111111111011011101011001100011001" & 
    "11111111111100100110100101100011011" & 
    "11111111111101000000101111000001001" & 
    "00000000000001000101100101011100000" & 
    "00000000000110011001110011001110100" & 
    "00000000001010100000001011010000110" & 
    "00000000001001110111010010000000110" & 
    "00000000000100010100101110110011011" & 
    "11111111111110111101101100001101011" & 
    "11111111111100010001000000000000111" & 
    "11111111111011100111100011010111010" & 
    "11111111111010101011000111111101010" & 
    "11111111111000101001110101011001001" & 
    "11111111110111000100001100110010000" & 
    "11111111111010001011111111011010101" & 
    "00000000000010001010010010011011111" & 
    "00000000001000111011011011011111100" & 
    "00000000001100110100110001011001111" & 
    "00000000001110010000001001110100010" & 
    "00000000001011001101110011010101101" & 
    "00000000000100100110111010011111011" & 
    "11111111111101010101100010011001000" & 
    "11111111111001100001100111111000111" & 
    "11111111111001101101010001110011001" & 
    "11111111111011110111100101111001100" & 
    "11111111111111010110010111011010010" & 
    "00000000000010010000010010001001100" & 
    "00000000000010101001111001011110101" & 
    "00000000000000110101001011000110011" & 
    "00000000000000011011011010110101110" & 
    "00000000000101100010010000010111100" & 
    "00000000001011111010101011101101011" & 
    "00000000001100011100010111100100011" & 
    "00000000000110111111000011111100111" & 
    "00000000000000000000101001010010001" & 
    "11111111111011100100110001011101111" & 
    "11111111111001011110000011010100001" & 
    "11111111110111100110001000100111111" & 
    "11111111110110010111101110010000001" & 
    "11111111110110101101011000001000011" & 
    "11111111111010011100000111011100110" & 
    "00000000000000000101001011101001010" & 
    "00000000000100111110110011000001000" & 
    "00000000000110111010011011000110101" & 
    "00000000000010101111010001000111000" & 
    "11111111111010000110111100011110011" & 
    "11111111110010010000101111001011111" & 
    "11111111110001011000100011001001001" & 
    "11111111110110110010010100011110001" & 
    "11111111111010100000011011001010011" & 
    "11111111111010001101101001011110010" & 
    "11111111111000110110101111010111101" & 
    "11111111111100001101010110011110111" & 
    "00000000000101000100010010001001111" & 
    "00000000001011111101001101101100001" & 
    "00000000001101011100011001111001000" & 
    "00000000001011100010101000010111101" & 
    "00000000001001000001101011011000101" & 
    "00000000000110000111111010011001101" & 
    "00000000000010110000011111100001001" & 
    "00000000000001011101111001000010110" & 
    "00000000000000011111111111011111110" & 
    "11111111111110110100011101001111001" & 
    "11111111111100101001111001101111001" & 
    "11111111111100001110101101001100011" & 
    "00000000000000110001110110111100101" & 
    "00000000000110111010110001110010111" & 
    "00000000001010100001111001111111100" & 
    "00000000001100000010010101001000110" & 
    "00000000001100011101001000100100101" & 
    "00000000001011000000111010010110000" & 
    "00000000000101000000101000111101000" & 
    "11111111111011001010110100100101111" & 
    "11111111110001100001001110111111011" & 
    "11111111101100010100010001010100111" & 
    "11111111101100001001001000010101100" & 
    "11111111101111110011011011011100010" & 
    "11111111111000111000001110000101010" & 
    "00000000000101010010110011010000110" & 
    "00000000001100101011101101100111101" & 
    "00000000001011010011111110001111010" & 
    "00000000000011101110110011100000000" & 
    "11111111111011011111111011000010111" & 
    "11111111110111111100110011001101101" & 
    "11111111111000000100101100100001000" & 
    "11111111111001011000110111000110001" & 
    "11111111111010101100100010100101101" & 
    "11111111111010100100001111010011001" & 
    "11111111111000000010000000100000101" & 
    "11111111110101111110100110000110100" & 
    "11111111111000100110000010010111110" & 
    "11111111111101110110110100011110111" & 
    "00000000000011110011010101011000101" & 
    "00000000001010000100100010101010110" & 
    "00000000001110001010011011011001010" & 
    "00000000001110011010101101001001001" & 
    "00000000001000001011110100000001100" & 
    "11111111111100110001010001111101000" & 
    "11111111110011011011001101010111011" & 
    "11111111110001110011110101010000100" & 
    "11111111110110101101010110111111000" & 
    "11111111111100000110000111001001011" & 
    "00000000000000100001101011101101010" & 
    "00000000000101000101001001000011000" & 
    "00000000001000001101001000010010001" & 
    "00000000001001000111000011010100001" & 
    "00000000000110100010001111110111111" & 
    "00000000000011100100010100101111001" & 
    "00000000000011000100001000110010000" & 
    "00000000000001001111100001101001000" & 
    "11111111111100000111110111100100101" & 
    "11111111110110100111100001100111001" & 
    "11111111110100110101110100111110001" & 
    "11111111111000100100100110110011010" & 
    "11111111111111001011011011000000101" & 
    "00000000000100111011000101010000011" & 
    "00000000000100100111010100011101110" & 
    "11111111111111100001000011000111011" & 
    "11111111111011000110100001101010110" & 
    "11111111111001100010111100011110010" & 
    "11111111111011101010000010001010101" & 
    "11111111111110001101110011101000000" & 
    "11111111111110101110011000001000111" & 
    "11111111111100111110111010011011010" & 
    "11111111111000100110111001001011111" & 
    "11111111110101110110111100010111111" & 
    "11111111110110110001000111001011000" & 
    "11111111111011000010100010101101011" & 
    "00000000000000011010001101010110011" & 
    "00000000000011111001001011001101001" & 
    "00000000000101101101000111001010011" & 
    "00000000000110101000111101101000110" & 
    "00000000000111000101111010010111011" & 
    "00000000000100101000010011100011100" & 
    "11111111111101011110000000010100000" & 
    "11111111110101110111111000011010000" & 
    "11111111110010000110011011100011101" & 
    "11111111110110010100001111001010111" & 
    "11111111111110101101000111101010001" & 
    "00000000000010111001010111011100110" & 
    "00000000000011011100110011100110100" & 
    "00000000000100010000011010011001100" & 
    "00000000000100111111001111101101111" & 
    "00000000000011110101111101100001010" & 
    "00000000000001000001110010001110110" & 
    "11111111111111010100000100101111010" & 
    "00000000000000110110101110111001111" & 
    "00000000000011000000100010100011011" & 
    "00000000000001100001000100110100110" & 
    "11111111111100010001010110100011010" & 
    "11111111111000010101001110000000011" & 
    "11111111111001011111101010000111110" & 
    "00000000000000100100000111010000011" & 
    "00000000001001111110000101001101010" & 
    "00000000001101110111110100111001111" & 
    "00000000001010011111111001101001011" & 
    "00000000000100111111111111001000100" & 
    "00000000000011101100010000100110100" & 
    "00000000001000110001000110000100010" & 
    "00000000001101110000011101110010000" & 
    "00000000001100101000011001000101101" & 
    "00000000000101100101000000110011010" & 
    "11111111111101101111011100110010001" & 
    "11111111111010100010001011111111011" & 
    "11111111111101001100111101000001100" & 
    "00000000000010100010110110101111101" & 
    "00000000000110101001011100010101101" & 
    "00000000001000000101001011111100001" & 
    "00000000000110101001101001001001110" & 
    "00000000000001110101100001101101001" & 
    "11111111111100110101001000001101001" & 
    "11111111111000100110101001000010111" & 
    "11111111110101011001110010111110101" & 
    "11111111110100001111101100001000010" & 
    "11111111110011001111000111110011001" & 
    "11111111110100011000000001111101111" & 
    "11111111111001010010010000111000000" & 
    "11111111111110111011100010001011110" & 
    "00000000000001010011101100010011110" & 
    "11111111111110111010010100111000111" & 
    "11111111111100010101001110011010100" & 
    "11111111111101000101010101001101010" & 
    "00000000000000010101011101110101110" & 
    "00000000000001111111011000110001011" & 
    "11111111111111100111111100101101101" & 
    "11111111111101100111001100001001100" & 
    "11111111111110010000111111000100011" & 
    "11111111111111000100000101011111100" & 
    "11111111111101010111011011011100110" & 
    "11111111111001111111011100000101001" & 
    "11111111111001111001101110011010101" & 
    "11111111111111100011100001001101110" & 
    "00000000001001010001100011100100001" & 
    "00000000010000011001001100000111000" & 
    "00000000001111101110011110110000010" & 
    "00000000001001001101111011001110111" & 
    "00000000000000101101001110000100100" & 
    "11111111111010000110111010111001110" & 
    "11111111110110000110100011001111110" & 
    "11111111110011100011100001101011100" & 
    "11111111110101010101011101110000010" & 
    "11111111111100100101101100010111100" & 
    "00000000000101011011001000110001100" & 
    "00000000001011001010101110011000110" & 
    "00000000001010111111001011111000110" & 
    "00000000000111010000010101111011000" & 
    "00000000000011011011001100001000001" & 
    "00000000000001100110000010111010100" & 
    "00000000000010010111001011011110110" & 
    "00000000000011101110101000001000110" & 
    "00000000000100000101101101100000001" & 
    "00000000000001111000010110010010101" & 
    "11111111111100100101111000001100111" & 
    "11111111110111010110101011101100001" & 
    "11111111110011101110111000101010101" & 
    "11111111110100010100011110100110011" & 
    "11111111111001111001101011111111000" & 
    "00000000000011010011101110110001100" & 
    "00000000001011110001010110110111111" & 
    "00000000001100100001001100111110001" & 
    "00000000000110100011110011101100111" & 
    "00000000000000110011101100110010000" & 
    "11111111111111110010111100010011111" & 
    "00000000000001110001011001111101010" & 
    "11111111111111101011101001100011101" & 
    "11111111111001111111110010001000010" & 
    "11111111110110010011111101001101001" & 
    "11111111111010100111001010011100110" & 
    "00000000000100001011001001000110001" & 
    "00000000001010101010000101001000000" & 
    "00000000001011010011001100100000000" & 
    "00000000000110101001110010110111010" & 
    "00000000000001000100000111100111111" & 
    "11111111111110101111010101100110000" & 
    "11111111111101101000001111000001000" & 
    "11111111111011110001010100100011011" & 
    "11111111111010010010100001001010000" & 
    "11111111111011111011001100111000111" & 
    "11111111111111101011101001011100111" & 
    "00000000000001100101001010111010100" & 
    "11111111111111101011100100001011100" & 
    "11111111111011110111000100011111110" & 
    "11111111111100011011101110011011100" & 
    "00000000000001011001000110010010101" & 
    "00000000000011110011010111011101100" & 
    "00000000000000110000001011101110110" & 
    "11111111111011011100011010010101110" & 
    "11111111111000010000010000011001000" & 
    "11111111111000100001101101111111001" & 
    "11111111111001001000110010000111011" & 
    "11111111111000001100110001001101111" & 
    "11111111110111000000111000101110100" & 
    "11111111111000110111100101111011011" & 
    "11111111111101001110111111000010110" & 
    "00000000000001101101100000000011111" & 
    "00000000000101010100011011011100000" & 
    "00000000001000110000111011101000111" & 
    "00000000001011001001101101001011000" & 
    "00000000001100000101100101101010010" & 
    "00000000000111111011011100010000101" & 
    "11111111111110111011111100100001001" & 
    "11111111110110010001110101001111011" & 
    "11111111110010111110010111111111001" & 
    "11111111110101111111011101011101110" & 
    "11111111111011111000111100111011111" & 
    "00000000000010101110111110010111111" & 
    "00000000001001000010010110011001011" & 
    "00000000001110001010100010100000101" & 
    "00000000010001000111000010001001010" & 
    "00000000001101100011100010101010010" & 
    "00000000000101010010010100001000010" & 
    "11111111111011100101010001011110011" & 
    "11111111110101101010000110010111110" & 
    "11111111110110010010001100001111010" & 
    "11111111110111110011111110000100000" & 
    "11111111111000110011101111111010011" & 
    "11111111111010110110111100101001110" & 
    "00000000000000100101001101110001100" & 
    "00000000001001110100011111111000001" & 
    "00000000010000110011111110010101001" & 
    "00000000010001111001000110111111110" & 
    "00000000001100111100100011000110100" & 
    "00000000000101011111000111100011111" & 
    "00000000000000010000100111101000011" & 
    "11111111111101100101001000001011011" & 
    "11111111111100011001010011000000010" & 
    "11111111111010111000110010000111000" & 
    "11111111111011010110000101101100101" & 
    "11111111111110001001001101011001001" & 
    "00000000000000001110110001010000111" & 
    "00000000000001001111100110001110111" & 
    "00000000000010011100111001100011011" & 
    "00000000000111011000011010001101100" & 
    "00000000001110001101110111000000110" & 
    "00000000001111000001101000101110001" & 
    "00000000001001111010011110001000100" & 
    "00000000000001110111011110010100111" & 
    "11111111111100000111101000101101101" & 
    "11111111111011000100010011010000011" & 
    "11111111111011010001000101111110101" & 
    "11111111111010100111110011000000100" & 
    "11111111111011101110000010101001001" & 
    "00000000000000101110001111101110110" & 
    "00000000000110011110011110011000101" & 
    "00000000001001100001101001110100111" & 
    "00000000001000010001101011000010001" & 
    "00000000000010010011011111010010110" & 
    "11111111111101111101110101101100100" & 
    "11111111111111101100100000111100110" & 
    "00000000000100001111101010011011000" & 
    "00000000000101101000101110001100111" & 
    "00000000000000100111001110010001111" & 
    "11111111111000111001100111000010011" & 
    "11111111110101111101010000010100111" & 
    "11111111111001110111111000000101111" & 
    "00000000000001010010011101001100100" & 
    "00000000000111101001000010100000000" & 
    "00000000001010001110010011001111011" & 
    "00000000000111110011010010010100001" & 
    "00000000000010011110010100000011110" & 
    "00000000000001001101010011111101000" & 
    "00000000000100111100100111000001110" & 
    "00000000000110001010100101011111100" & 
    "00000000000000111101100100100101001" & 
    "11111111110111111101111110011001111" & 
    "11111111110010110101100001100110101" & 
    "11111111110111001111010001010011011" & 
    "00000000000010110101010000010100000" & 
    "00000000001101111000111001100010000" & 
    "00000000010010000000010011000000010" & 
    "00000000001111101000101100001110010" & 
    "00000000001010010101101101011011111" & 
    "00000000000110011001011101011000111" & 
    "00000000000101001011000010110010110" & 
    "00000000000100010010101101000001100" & 
    "00000000000011001011110110110000010" & 
    "00000000000000001001011101111001110" & 
    "11111111111100111001001100111110101" & 
    "11111111111100101010000000011111111" & 
    "11111111111101110110111101100001101" & 
    "00000000000001101010000100110010000" & 
    "00000000000110111001100110000001011" & 
    "00000000001011001111110011100001010" & 
    "00000000001101101110111010111110011" & 
    "00000000001100111101011010010100101" & 
    "00000000001011110111000010101110111" & 
    "00000000001010000111001000011101101" & 
    "00000000000011101101111111001110100" & 
    "11111111110111111110001000111011000" & 
    "11111111101101010100100000010110011" & 
    "11111111101101100100101101001101000" & 
    "11111111111000011101101010101110011" & 
    "00000000000110100000010011000111001" & 
    "00000000010000010111001011001010000" & 
    "00000000010001011011100010100111101" & 
    "00000000001100011000100000110101001" & 
    "00000000000111000111100000010100011" & 
    "00000000000101000011001110001011100" & 
    "00000000000011101001011100001001001" & 
    "11111111111110110110110000011010110" & 
    "11111111111000101111111010001000000" & 
    "11111111110101010001100001000110010" & 
    "11111111110110111100001000101001011" & 
    "11111111111010111111010000000010111" & 
    "11111111111011110000111100010010000" & 
    "11111111111011000010100001101111000" & 
    "11111111111010100010011001100001011" & 
    "11111111111100110111000111100001111" & 
    "00000000000010010110011101011110110" & 
    "00000000000101101010101111110000001" & 
    "00000000000010011001010001011001110" & 
    "11111111111010110010011110011011011" & 
    "11111111110101011010110011100010101" & 
    "11111111110110000110000100000111000" & 
    "11111111111010001001001110010101011" & 
    "11111111111111010010101001011110010" & 
    "00000000000010010011010100110110011" & 
    "00000000000010101101011000001101111" & 
    "00000000000100111001011010110100101" & 
    "00000000001001010001000111010100100" & 
    "00000000001100010101101000011101010" & 
    "00000000001010001011000001010101110" & 
    "00000000000011001000011010001000100" & 
    "11111111111100011101000000011100110" & 
    "11111111111000100100001100110111111" & 
    "11111111110111100110001101000110110" & 
    "11111111110111000101001010110000011" & 
    "11111111111001000010000101111101110" & 
    "11111111111100111010000001011101010" & 
    "11111111111110010111001010100111101" & 
    "11111111111111000010001101010100110" & 
    "00000000000000010000001101101101110" & 
    "00000000000010001010010110101111100" & 
    "00000000000011001101101011011001110" & 
    "00000000000001110111010100001010000" & 
    "00000000000000010010010100001011110" & 
    "11111111111111011001110010111111110" & 
    "11111111111111101001000111111001000" & 
    "00000000000000011100010101010010111" & 
    "11111111111111011011100100000011011" & 
    "11111111111011100111010100110001010" & 
    "11111111110111010010000110000111001" & 
    "11111111111001001110101011110101100" & 
    "00000000000011010100010111011100111" & 
    "00000000001110010001011011100010100" & 
    "00000000010001000010110011001011100" & 
    "00000000001001101000000111100011001" & 
    "00000000000000110111000000000011011" & 
    "11111111111101001001110111110010001" & 
    "11111111111100011101111111011001011" & 
    "11111111111001101110011110111001110" & 
    "11111111110011100110111000110100111" & 
    "11111111101110101101101000111110000" & 
    "11111111110001101011001011111000001" & 
    "11111111111010100110011111010011101" & 
    "00000000000011011001011101100110110" & 
    "00000000001000010110101111011001010" & 
    "00000000001001010111011011101101101" & 
    "00000000001000111011011111100001100" & 
    "00000000001001000001000010111001010" & 
    "00000000001000011001110110011111010" & 
    "00000000000101011001011101111000110" & 
    "00000000000000111010011001110011000" & 
    "11111111111100001110101011100111101" & 
    "11111111110101111100101010001100010" & 
    "11111111110010100001010110010001100" & 
    "11111111110011111110100111011111111" & 
    "11111111111001001101101110010100100" & 
    "00000000000000011100011110101000001" & 
    "00000000000101110111111000110001110" & 
    "00000000001001011100001111001101001" & 
    "00000000001010110101000101110000001" & 
    "00000000001000010011101111111011011" & 
    "00000000000010110011010011001000100" & 
    "11111111111101110110111100111100000" & 
    "11111111111100011000011110111001110" & 
    "11111111111010101101000101011101001" & 
    "11111111110111110010100000000101001" & 
    "11111111110111100011001001100100001" & 
    "11111111111101011101010000111000101" & 
    "00000000000110101111101111011010100" & 
    "00000000001001111101001011011111000" & 
    "00000000000100111001110110101111101" & 
    "11111111111110111000100010100111100" & 
    "11111111111111000010110010100001011" & 
    "00000000000010111001010111110101011" & 
    "00000000000011110100001101101001000" & 
    "00000000000000101010101000010100010" & 
    "11111111111110001011010000000001010" & 
    "11111111111110100110100010111011001" & 
    "11111111111111000111110010011110101" & 
    "11111111111100100100010100101001010" & 
    "11111111111010001000011100011111011" & 
    "11111111111110101110101011110011111" & 
    "00000000001001100101010001000000010" & 
    "00000000010001010111101100111011110" & 
    "00000000001111000111011110011101010" & 
    "00000000000110101100010110110101001" & 
    "00000000000000111111110111110011111" & 
    "11111111111110101101101110101011110" & 
    "11111111111010111110111001101100000" & 
    "11111111110100001000101000001101000" & 
    "11111111110000101101110011011010000" & 
    "11111111110110011100000001011100101" & 
    "00000000000000010011011010111110000" & 
    "00000000000110101001110001111000001" & 
    "00000000000111101100010100010000000" & 
    "00000000000111010000110000010111110" & 
    "00000000001000101000010010110000110" & 
    "00000000001001011011010110011111100" & 
    "00000000000111010010100101111000100" & 
    "00000000000001001010111101101011010" & 
    "11111111111001000111100010111010001" & 
    "11111111110011110100111111111111111" & 
    "11111111110100110101000111000011111" & 
    "11111111111101010111100000000111110" & 
    "00000000000111100100110000010111010" & 
    "00000000001100010011000100111111101" & 
    "00000000001010001111010101001100010" & 
    "00000000000101011000110000110011100" & 
    "00000000000011001001010110110110110" & 
    "00000000000010000011111101011001100" & 
    "00000000000000001100001101101101111" & 
    "11111111111101001111100010011101111" & 
    "11111111111001100101111110100110110" & 
    "11111111110110111011000110100010111" & 
    "11111111110110110011101001111001010" & 
    "11111111111010001010110000111110100" & 
    "11111111111110011010010110000011001" & 
    "00000000000001110010011100100110001" & 
    "00000000000110000111000000001011010" & 
    "00000000001010010010101101110101000" & 
    "00000000001110001101101110010100001" & 
    "00000000001111011110110011110001111" & 
    "00000000001001110011011101000011111" & 
    "00000000000001001111000010100001000" & 
    "11111111111100001001011010111010000" & 
    "11111111111100001010000101011011011" & 
    "11111111111100111010110101101000111" & 
    "11111111111010101001010011011001101" & 
    "11111111110110101100000110010011110" & 
    "11111111110100011110101101100000001" & 
    "11111111110110111100011011000011101" & 
    "11111111111011011100110101011100111" & 
    "00000000000000101001000011101010001" & 
    "00000000000111001110001011101100001" & 
    "00000000001100000001110101101001111" & 
    "00000000001011011010100000010110010" & 
    "00000000000110010001110111111011110" & 
    "11111111111110100101111011101011101" & 
    "11111111110110110110011000001101110" & 
    "11111111110010000101101111100110010" & 
    "11111111110010111110001100001011000" & 
    "11111111111000010110001010100110100" & 
    "11111111111101010110110100011110010" & 
    "00000000000010011010101110110101110" & 
    "00000000000111110111101101001111011" & 
    "00000000001010111011110001111001011" & 
    "00000000000111011100111110111011100" & 
    "11111111111101001101100111110101101" & 
    "11111111110101111111101110011000000" & 
    "11111111110101111011010101100001101" & 
    "11111111111010000001100001110010010" & 
    "11111111111101010101010010111111001" & 
    "11111111111101100010100000101010101" & 
    "11111111111100101001100101000011100" & 
    "11111111111001101011010111110001001" & 
    "11111111110110101100000111011111001" & 
    "11111111111000110101000101101101010" & 
    "00000000000000010101100010001100100" & 
    "00000000000111001101000101101000111" & 
    "00000000000110001011101000010001011" & 
    "11111111111111111001111101111110101" & 
    "11111111111011100101100111001001010" & 
    "11111111111011010100011111100101000" & 
    "11111111111101001001000001001101011" & 
    "11111111111101100010010100000001101" & 
    "11111111111100001100010000000000011" & 
    "11111111111011000010010001111110100" & 
    "11111111111011110101110110100011111" & 
    "11111111111111010001110001111011101" & 
    "00000000000001011110101010000101111" & 
    "00000000000001000101001000001011010" & 
    "00000000000001111000011000000111100" & 
    "00000000000100100110000111000100111" & 
    "00000000000110000111010001001000000" & 
    "00000000000010001101110100010100000" & 
    "11111111111010000010110110000111100" & 
    "11111111110100011111010100001010101" & 
    "11111111110100110000011011000001111" & 
    "11111111111001011110000001101100001" & 
    "11111111111101001110111101010001011" & 
    "11111111111111001010010011100000100" & 
    "00000000000001110100000010110010010" & 
    "00000000000101110010011101011000010" & 
    "00000000001010110101010110111001110" & 
    "00000000001101011111011011110001100" & 
    "00000000001011000011101010111101100" & 
    "00000000000100011101111101110000110" & 
    "11111111111101010111111011011000110" & 
    "11111111111010100000101100100000111" & 
    "11111111111001101110001011000100010" & 
    "11111111111001100011100111101110011" & 
    "11111111111011000101010100110101001" & 
    "11111111111110101011110110010011101" & 
    "00000000000100001000001001001010010" & 
    "00000000000111111001111001111100111" & 
    "00000000000111111001100100110000110" & 
    "00000000000110111010110001010110111" & 
    "00000000000110011011001001000100100" & 
    "00000000000110011011011001001101101" & 
    "00000000000100011010010101111100000" & 
    "00000000000000110000100101111100110" & 
    "11111111111011100001001010101010011" & 
    "11111111110100000011110010001010100" & 
    "11111111101111001111100101000000111" & 
    "11111111110011001000100011110010101" & 
    "11111111111111010110001010111001011" & 
    "00000000001011001001110111010010111" & 
    "00000000001110010100011010101110110" & 
    "00000000001011010111011010110011001" & 
    "00000000000111101010101001000100100" & 
    "00000000000111101110000100011011011" & 
    "00000000001001011000010100110101011" & 
    "00000000000110100001110101101001000" & 
    "11111111111101111101101111110010101" & 
    "11111111110011010011011000011101011" & 
    "11111111101101100100011101010101100" & 
    "11111111101111011110000000111110111" & 
    "11111111110110111100111111010100000" & 
    "11111111111111110100101110011100011" & 
    "00000000000101001101000010110011101" & 
    "00000000000110110000101011010111010" & 
    "00000000000101001011111001101010111" & 
    "00000000000000110000011001100001111" & 
    "11111111111101011100010000101011111" & 
    "11111111111100010100010000100101110" & 
    "11111111111010010111000010110101100" & 
    "11111111110110001001100111111010111" & 
    "11111111110011100001100101110101110" & 
    "11111111110100101101000010000111011" & 
    "11111111111001010000110111000110110" & 
    "11111111111110111001101101110111110" & 
    "00000000000011001100110100011000011" & 
    "00000000000101101000101110010000111" & 
    "00000000001001101010101111101001110" & 
    "00000000001101101010001110110110011" & 
    "00000000001101101001110000100010111" & 
    "00000000001001000101010100011110100" & 
    "00000000000000100011111110111000010" & 
    "11111111111000000101110100100101011" & 
    "11111111110100100100101000100011001" & 
    "11111111110101101010010110110001110" & 
    "11111111111000001001000111001011011" & 
    "11111111111011011110100010111101101" & 
    "00000000000010010011000101110110000" & 
    "00000000001010110111110110011001011" & 
    "00000000010001010010100010111101110" & 
    "00000000010001011000000110111000011" & 
    "00000000001001111011011001010110101" & 
    "00000000000001101000110011000110010" & 
    "11111111111101100110010110010100110" & 
    "11111111111011001001100011001101011" & 
    "11111111110111000110001101011101100" & 
    "11111111110001111101110001011110100" & 
    "11111111110000001001001111111100101" & 
    "11111111110100001111101110101111001" & 
    "11111111111100000100100101101011110" & 
    "00000000000100110011010011010000101" & 
    "00000000001011011110100000000100011" & 
    "00000000001101101100000010010111110" & 
    "00000000001000110010110100001011100" & 
    "00000000000000110101001010110001101" & 
    "11111111111011101110001100110000000" & 
    "11111111111010001010001000100000010" & 
    "11111111111010101101000100010110100" & 
    "11111111111010001101111011110000011" & 
    "11111111111001011110000111001011010" & 
    "11111111111010101101000111100000100" & 
    "11111111111110000111101001110000100" & 
    "00000000000101000101101011001010001" & 
    "00000000001011101000010110010011111" & 
    "00000000001100110011011010000110000" & 
    "00000000001000000100010110111110111" & 
    "00000000000010100111110101011001100" & 
    "00000000000000100010111111111000110" & 
    "00000000000000101000100110110111000" & 
    "00000000000000010001100110000010000" & 
    "11111111111101010100011110100001101" & 
    "11111111111001001111110101100000100" & 
    "11111111110110100101000011110100110" & 
    "11111111110110011000010111111010100" & 
    "11111111111010100011101100010010110" & 
    "00000000000001110110000001000000100" & 
    "00000000000111000001010101111100010" & 
    "00000000001001000101100110100010010" & 
    "00000000001010010100101000001110000" & 
    "00000000001010011110100110111010010" & 
    "00000000001000001111010000010110010" & 
    "00000000000001100100100101111111110" & 
    "11111111110111001101011001010101001" & 
    "11111111101111110110000010110100000" & 
    "11111111110001100001011011011111101" & 
    "11111111111001100001111111110100101" & 
    "11111111111111100000100011000010110" & 
    "00000000000010001111011100111001001" & 
    "00000000000010110001010111110101100" & 
    "00000000000100011110100101100110101" & 
    "00000000000111001001100110100101010" & 
    "00000000000110110001011011001001011" & 
    "00000000000010000011011100001000110" & 
    "11111111111010101010111100111001111" & 
    "11111111110101000001010110001011100" & 
    "11111111110100000000111001011101001" & 
    "11111111110110001111100101011111010" & 
    "11111111111001010001001001011000010" & 
    "11111111111011011101101000100010011" & 
    "11111111111111000010001001101010001" & 
    "00000000000101011010101100100110111" & 
    "00000000001100000101000110001010110" & 
    "00000000001110110001010111001101111" & 
    "00000000001100000111000010001101101" & 
    "00000000000101110000011001010010010" & 
    "11111111111111100001001111100011001" & 
    "11111111111100001101001101011110011" & 
    "11111111111011110000010010101101000" & 
    "11111111111001111101100110101110010" & 
    "11111111110110110110010110100100100" & 
    "11111111110111100010100011001101001" & 
    "11111111111011110101011100110100001" & 
    "00000000000001011011110000010101001" & 
    "00000000000101100111010110000011010" & 
    "00000000001000010011110110111100101" & 
    "00000000001010101111011101000110001" & 
    "00000000001001001001100101001011111" & 
    "00000000000010001100110101011000110" & 
    "11111111111001011000111010111101001" & 
    "11111111110101010100101000111101100" & 
    "11111111110101100000010001111000011" & 
    "11111111110101011100110111000110010" & 
    "11111111110111001010110100001101110" & 
    "11111111111010101111001001010011100" & 
    "11111111111111100000010011001000110" & 
    "00000000000011110010100101010000101" & 
    "00000000000101011111011100001010011" & 
    "00000000000111001100111010100111110" & 
    "00000000001001111001011100001000011" & 
    "00000000001000101011000101000101000" & 
    "00000000000000000111000010010110110" & 
    "11111111110101100110111110101111110" & 
    "11111111110000000101111110011101000" & 
    "11111111110000111101100001000101100" & 
    "11111111110101010010110101010010111" & 
    "11111111111000110110111011110101000" & 
    "11111111111011111101100011001100010" & 
    "00000000000000110111011101110000010" & 
    "00000000000101000110111001110100100" & 
    "00000000000110011011110010111110011" & 
    "00000000001000001111010100010011010" & 
    "00000000001010101001000000011101010" & 
    "00000000001010011010111001100100011" & 
    "00000000000011110110110001100111010" & 
    "11111111111001101001001111111000010" & 
    "11111111110100100001001000101001000" & 
    "11111111110110111110000110110001101" & 
    "11111111111100011111100011100010010" & 
    "11111111111110110000011000101100000" & 
    "11111111111111000110100010010010000" & 
    "00000000000011111101110111101010010" & 
    "00000000001100100011111011101010110" & 
    "00000000010010100100010001000001001" & 
    "00000000010000100010010110001011001" & 
    "00000000001000011101110111100111110" & 
    "00000000000000011110110010001111011" & 
    "11111111111011010010110000100111000" & 
    "11111111111001100011001010010000011" & 
    "11111111111001101011101101011001001" & 
    "11111111111011001111011010110001101" & 
    "00000000000000010100010101000001000" & 
    "00000000000111010110011011111101011" & 
    "00000000001011101011101011110010100" & 
    "00000000001001100110011100100100100" & 
    "00000000000001111111111011010001011" & 
    "11111111111010111000000101111000001" & 
    "11111111111000001001100010011110110" & 
    "11111111111001100101011101000101100" & 
    "11111111111011010010101011010111100" & 
    "11111111111100000001111101001110110" & 
    "11111111111011000101100111001101110" & 
    "11111111110111011011110111010101000" & 
    "11111111110110001001000100011111010" & 
    "11111111111000110011010000010101101" & 
    "11111111111100100101011000110011110" & 
    "11111111111111111101001111001010001" & 
    "00000000000001111000000111100100000" & 
    "00000000000100011110100101010110110" & 
    "00000000000111100010111110101111100" & 
    "00000000001000001100111001110101100" & 
    "00000000000101000000001110110001001" & 
    "11111111111111101110001000011110111" & 
    "11111111111011110000110010111101010" & 
    "11111111111000110110011101100010101" & 
    "11111111110110101010101100011101000" & 
    "11111111110101110001111111110011000" & 
    "11111111110111010011011001010101010" & 
    "11111111111101110000100010001110111" & 
    "00000000000101011101100100000100011" & 
    "00000000001001101001000000001010110" & 
    "00000000001001011010001110100100000" & 
    "00000000000111000010010001101101001" & 
    "00000000000101011001001010011101001" & 
    "00000000000011001011101101001001001" & 
    "11111111111111100101001000010101111" & 
    "11111111111011100000000001010111010" & 
    "11111111110111101000100101110011001" & 
    "11111111110100001111011000101011111" & 
    "11111111110011000011101100110010011" & 
    "11111111110111001010000100101000101" & 
    "00000000000000010100001111011000100" & 
    "00000000001001000001100001111000010" & 
    "00000000001101011111100111000111001" & 
    "00000000001110111001001001011110101" & 
    "00000000001110111001000110000110000" & 
    "00000000001011010001000111010101101" & 
    "00000000000001111000011010110010000" & 
    "11111111110111100000001110011000110" & 
    "11111111110100000101001111101011110" & 
    "11111111111010001101100110100000111" & 
    "00000000000010110010101001000101011"
  );

end pkg_OutputSamplesFi;
