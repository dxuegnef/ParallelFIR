
library ieee;
use     ieee.std_logic_1164.all;


package pkg_InputSamplesFi is

  type T_INPUTSAMPLESFI is array (0 to 2501-1) of std_logic_vector(16-1 downto 0);

  constant PKG_INPUTSAMPLESFI : T_INPUTSAMPLESFI := (
    "0010100010011010",
    "0001111001101011",
    "1110100101100000",
    "0001001110111110",
    "1111000101011000",
    "1110111000100010",
    "1101110000111111",
    "1111101110001101",
    "0011010000000000",
    "0001110001011110",
    "1111111101011001",
    "0010111101000111",
    "0010000000001100",
    "0001001101101111",
    "0000101000101000",
    "0001000110101010",
    "1110111000010010",
    "0001001010010101",
    "0000110010011101",
    "1111100111011011",
    "0000110111001101",
    "1101100011101100",
    "0001000101101101",
    "0010011110011010",
    "0000100011100110",
    "0011000010001110",
    "0000110010110101",
    "0000100010101010",
    "0000101010100111",
    "1101111110100110",
    "0001000101000101",
    "1101000011010100",
    "1110010011110111",
    "1110110111001011",
    "1100000011110011",
    "0010101111110101",
    "0000001111101100",
    "0000100001011101",
    "0010101001011110",
    "1110001101010110",
    "0001001101001111",
    "1110110000110010",
    "1111111111011010",
    "1111101100010011",
    "1101010101011000",
    "0000001010010011",
    "1110100110011011",
    "0000111111111110",
    "0001111100000010",
    "0001001011010011",
    "0001001000101110",
    "0000001001010000",
    "1111101000010111",
    "1111010000100010",
    "1110110000100010",
    "0001101110010100",
    "1101011011011110",
    "1111110000000011",
    "1111011100100011",
    "0000000111101111",
    "0000001110000101",
    "1111111100111101",
    "0001110101001000",
    "0010011000001101",
    "0001011101101101",
    "0001011001010010",
    "1101100000110001",
    "1110111011011110",
    "1110010100010101",
    "0000100011001010",
    "1111100100110101",
    "1111100000110110",
    "0000001011011111",
    "0001101110111100",
    "1111010011010111",
    "0000100110010000",
    "1110101001010010",
    "0001010101010100",
    "0000001100011100",
    "1110100100011011",
    "0001100111000100",
    "1110011111011001",
    "1111100100111100",
    "0001010000100110",
    "1110001100110000",
    "0010000000010111",
    "0000110000010101",
    "0001000010001011",
    "0001011111100100",
    "1110110000010001",
    "0000001010010100",
    "1111000110111100",
    "0000011001001101",
    "0001111101110000",
    "1101100010000011",
    "0000011000001110",
    "1110101011101100",
    "1110011100000101",
    "0000011001111110",
    "1110010001011101",
    "0010110101110010",
    "1111001011011110",
    "0000111100011110",
    "1111110100111101",
    "1111000100011001",
    "1111100101110011",
    "1110101100000101",
    "0000000111100110",
    "0001011000100011",
    "1110110011110100",
    "1111001010111011",
    "1111000101001001",
    "0010101000011101",
    "0000001101001010",
    "0000111000011000",
    "0001011011101110",
    "0000011100001011",
    "1101101101011111",
    "1111001011101000",
    "1100111111011011",
    "0011000110010101",
    "1111100101110010",
    "0001110000000011",
    "1111110010010110",
    "1111100110010100",
    "0001101110100100",
    "0001001010100111",
    "0000100100010010",
    "0001000100101100",
    "1100101101101010",
    "1111110101100101",
    "1101011000000001",
    "1101110011010110",
    "0000001011100000",
    "1111010010010010",
    "0001010101111011",
    "1110100101100001",
    "0010011001111011",
    "0001101000001011",
    "1111100111101111",
    "0001010101001111",
    "1110101111011110",
    "1101111010111110",
    "1111000101111111",
    "1101010111100001",
    "1111001101100011",
    "1101100110111110",
    "1111110101101001",
    "1110110101111010",
    "0001000010000001",
    "0010100001010010",
    "0000000011000010",
    "0000110011110110",
    "1111100100101110",
    "1111110010001011",
    "0000000011101101",
    "1101011111000000",
    "0000101110110001",
    "1111011100100110",
    "1110011010100010",
    "0001000000111111",
    "1111000100100111",
    "0000001010000101",
    "0011110011011100",
    "0001100100110101",
    "0001100111011101",
    "1101101111110010",
    "1110110011100110",
    "1111001100111110",
    "1110111111011000",
    "1110110110111110",
    "1100011011110111",
    "1110111011000011",
    "0001001011011011",
    "0000011101010111",
    "0010011100111010",
    "1111111011111110",
    "0001000001110101",
    "1111111001010101",
    "1111101000001001",
    "1110110101000101",
    "1110101001110110",
    "1110100001111101",
    "1111010101100011",
    "1111100011100111",
    "0010010110010010",
    "1110110011010110",
    "0010100010011101",
    "0001111100000001",
    "1111110110100010",
    "0001000111010010",
    "1110110010010011",
    "1111010111100101",
    "1111011001110000",
    "1110010000000001",
    "0001000001000110",
    "0000010010101101",
    "0000110101101011",
    "0000101000101001",
    "0000101100010100",
    "0010001011101110",
    "1111000010011010",
    "0001110010110100",
    "0000101011011101",
    "1110111001101000",
    "0000101101001101",
    "1110011101011101",
    "1110011100000001",
    "1111100000100110",
    "1110110110111001",
    "0000110001101111",
    "0001100110100010",
    "0000011001101110",
    "0000110010110011",
    "1111001101010100",
    "0000001000101000",
    "1110110011111011",
    "1111011001011100",
    "0000111010001101",
    "1101111100110011",
    "1111001000000111",
    "0000010111100110",
    "0001100110110100",
    "0000100111011000",
    "1110100011111010",
    "0001100011100011",
    "1111111010010101",
    "0001000111101111",
    "0000000111000101",
    "1111001101010111",
    "0000100101010011",
    "1100111100101100",
    "1110011011100111",
    "1110111011100011",
    "1110011111101111",
    "0000111111010001",
    "1111111011101011",
    "1110001111111010",
    "0000110100100001",
    "0001001010011001",
    "0000001111100001",
    "1111111011111111",
    "0000000001011010",
    "1111010110011011",
    "1110011000011010",
    "1110101000000100",
    "1110101011100100",
    "0001111110011101",
    "0000111100010111",
    "0000000110111101",
    "0001010001000001",
    "0000000010010101",
    "0001000100111100",
    "0000110011000101",
    "1110011001000111",
    "1111111101000110",
    "0000001110010000",
    "1101000111101111",
    "0001111001101011",
    "1111010101110101",
    "0010010011110010",
    "1110010000011000",
    "0000101100000000",
    "0000111111111110",
    "0000010101111100",
    "1111101000111001",
    "1111011110011011",
    "1110011101010111",
    "1111011100100000",
    "1110110110011111",
    "0000100001001010",
    "1111110110010001",
    "0001011000001100",
    "0000001100011010",
    "0000010100110001",
    "0001000011100100",
    "1110101111101110",
    "0001110001010001",
    "0000010111110011",
    "1110101101011101",
    "0001000110100010",
    "1110110010110010",
    "1111101110101100",
    "0000111011000000",
    "1111111011101111",
    "0001100011001000",
    "1111001110101100",
    "0000101000000100",
    "0010011110000100",
    "1110010011101110",
    "0001010010001110",
    "1101000011100000",
    "0000101100010011",
    "0000001111011011",
    "1110001100110011",
    "0000000111101100",
    "1100010001110110",
    "0000111100111111",
    "1110101001110000",
    "1101101111111000",
    "0010000101000111",
    "1111000111100111",
    "0001010000011010",
    "0001000011001000",
    "1111100111111000",
    "1111011111111111",
    "1110101001011111",
    "1111011110101110",
    "0000011111110110",
    "1111100010100011",
    "0010001101001111",
    "1111110010011100",
    "0001001000010110",
    "0010010010010001",
    "1101110010111110",
    "0000110011011111",
    "1101101110111010",
    "1111010010100000",
    "0000000001110010",
    "1111000001100101",
    "1111001011010001",
    "1110010010110101",
    "0000100000100100",
    "0000100011011001",
    "0000010111101000",
    "0010011001100110",
    "1111001000110010",
    "0000101010110000",
    "1110001111010110",
    "1111111010010010",
    "1111100011111110",
    "1100111111101100",
    "1111001000000001",
    "1110001111100011",
    "1110111110111001",
    "0000101111111001",
    "0010000110010000",
    "0010011010101000",
    "1110110001111110",
    "0000010111001000",
    "1111111010010011",
    "1110101111111010",
    "1111110101100000",
    "0000001000001000",
    "1101111011010000",
    "0001110001000111",
    "1110010010001100",
    "0000101100110000",
    "0001100000100111",
    "0000001001110001",
    "0010111000011000",
    "0000011000111111",
    "0000000011111001",
    "1110100100010000",
    "0000100111111011",
    "1111100101100010",
    "1110010011010110",
    "1111111100010100",
    "1111110010010000",
    "1110000110010101",
    "0000110101110110",
    "1111110010111001",
    "0010110000011011",
    "0000011010101011",
    "0000101101000110",
    "0001100111100010",
    "1110110001010001",
    "1110100111010101",
    "1111000110000110",
    "1110000111001011",
    "1110101110001100",
    "1110111101010001",
    "1111100011001011",
    "0000110000000010",
    "0000011001110101",
    "0001000110000111",
    "1111110001110111",
    "0001001100011110",
    "1110100010010011",
    "1111110011010010",
    "0010100111011001",
    "1111001010001000",
    "1111000100000100",
    "0000000110011010",
    "1101111101111011",
    "0011001011111101",
    "0000110111000101",
    "0010000100001010",
    "0000011001101101",
    "0000001111010111",
    "0000110000000011",
    "1110101100010011",
    "1111000110100000",
    "1110010110101000",
    "1101010010100100",
    "1111111110110011",
    "1101000100010000",
    "0000111110101100",
    "0000101110100010",
    "0000110001000011",
    "0010010001010000",
    "0000100011111100",
    "1111010111001010",
    "1111010110100000",
    "1110010100010111",
    "0000010011001111",
    "1111010100111110",
    "1111000101101110",
    "0000111011101110",
    "1111011110101010",
    "0010011110111011",
    "0000000011000000",
    "0000100111101111",
    "1111110010111101",
    "0000000100110101",
    "0010001000001011",
    "1110101101100000",
    "1111001000011000",
    "1111000100100001",
    "1101000110100011",
    "1111101100101011",
    "1110100101011010",
    "0000011010101111",
    "0000110001111111",
    "0000101011011100",
    "0010000111000000",
    "0001111000011010",
    "0001001010000011",
    "0010001011010010",
    "1110000010101100",
    "0000101101111011",
    "1101111100000101",
    "1111111110101100",
    "0000010001000000",
    "1100110100010101",
    "1111111110110110",
    "1110011110101010",
    "0001101011011111",
    "0010101111110111",
    "1111100101111101",
    "0010000111110001",
    "1111100011001001",
    "1110100111101011",
    "1111110001101101",
    "1101011100100111",
    "0001101101010001",
    "1110101110111001",
    "0010000000100000",
    "0000011010110111",
    "0000101010000010",
    "0001111011111111",
    "1110000010111010",
    "1111110111001110",
    "0000111111000000",
    "1110101101011101",
    "1111000100101000",
    "1101100100101001",
    "1111101000001111",
    "1110101011011011",
    "1111111110101000",
    "0000101010110001",
    "0001101110101001",
    "0000001100101010",
    "0001011110100001",
    "1110011001100010",
    "0000100101011110",
    "1110011010010001",
    "0000000100101011",
    "0000010100100100",
    "1110011111111101",
    "1111110100010110",
    "1111100101001011",
    "0001001010111011",
    "0000111101110001",
    "0000101000110111",
    "0010011010011011",
    "1111000101001001",
    "0001100110101100",
    "1111101101101111",
    "1110001010010101",
    "0000010111100011",
    "1101111001000011",
    "1111001111110101",
    "0000010001000101",
    "0000000011001111",
    "0001000111000111",
    "0000001111110110",
    "0001000010100001",
    "0001100000011101",
    "0000010111000010",
    "0000101100010011",
    "1111010001110100",
    "0000010001011101",
    "1111011110001011",
    "1111111011011100",
    "1111100101010010",
    "1110000001110011",
    "1110100111110011",
    "0001110000010110",
    "0000111011110011",
    "0001111010111001",
    "0000111101110100",
    "0001000001110101",
    "0000101010011010",
    "1110111000001101",
    "0000101000011000",
    "1110010011001111",
    "0010001010101010",
    "1110100000010100",
    "1101001001100100",
    "0000001010110010",
    "1110110100111010",
    "0000110110000001",
    "0001000110111111",
    "1111101100111001",
    "0001110110011011",
    "1111011001001001",
    "0000011011000100",
    "0001001010000101",
    "1111011011000000",
    "1110111010000110",
    "1100011011111011",
    "0001010001100001",
    "1111000000100110",
    "0000001000100101",
    "0010000010010001",
    "0010010010110110",
    "0000110001101001",
    "1111110111010101",
    "1111000000000100",
    "0000011011111101",
    "1110010001001101",
    "1110110001010101",
    "1110011100101111",
    "1111010100011111",
    "1111111101110101",
    "1110111000110100",
    "0010100110111110",
    "0000110110111101",
    "1111110001111001",
    "0010001101010111",
    "1110101101000001",
    "0000101100110111",
    "1111000010001100",
    "1111001101100011",
    "0000110100100000",
    "1110100011010110",
    "1111100000011001",
    "1111110011010100",
    "1111110011000001",
    "0001100011111101",
    "1111101010001010",
    "0001110101000001",
    "0000000100110000",
    "1111111010001011",
    "1111101010001101",
    "1111001010111110",
    "1110110110110110",
    "1111110110010010",
    "1111111110010111",
    "0000111001010010",
    "1111011110110101",
    "0011010001111111",
    "0010001110101000",
    "1111011111001111",
    "0001111101010100",
    "1110101001001100",
    "0000011000001010",
    "0000110010111001",
    "1100100110000010",
    "0001001110000100",
    "0000001110010010",
    "0000011010110101",
    "0010100101110101",
    "0000001110010000",
    "0000110000110101",
    "1101110111111011",
    "0000100000101111",
    "0001000101011110",
    "1111000101010010",
    "0000100110101100",
    "1101100111110011",
    "1111100001011111",
    "1110000010000111",
    "1110001111100101",
    "0000011111011000",
    "0000011100001001",
    "0001010000110111",
    "0000000111110100",
    "1111111010010001",
    "0000100111101000",
    "1110010101100100",
    "0000100010010010",
    "1111011111100010",
    "1110100110001110",
    "0001000100110011",
    "1110111100100001",
    "0000111011000011",
    "0001100001110010",
    "0001001111001110",
    "0010011110011101",
    "0001011110101100",
    "0000110111100001",
    "0000010100101111",
    "0000011101110111",
    "1111101011100110",
    "1110001100100011",
    "0000010011001001",
    "1111110100100100",
    "0000011010001001",
    "0010010101111101",
    "0000001101100010",
    "0000100000000000",
    "0001110110000010",
    "1110100010011001",
    "0001100011011011",
    "1111110011111110",
    "1111111000100111",
    "0000010000100101",
    "0000001111001110",
    "0001000111010111",
    "1111000010000100",
    "0001000000110111",
    "0001010001010011",
    "1110110000001011",
    "0001100101010110",
    "0001010010101100",
    "0000110011010010",
    "0000111101000101",
    "1101110000100100",
    "0000010000010111",
    "1110110011001001",
    "1110000001001001",
    "0000000001001111",
    "1110110100100110",
    "0000010111101001",
    "1111111000011110",
    "1111011000011010",
    "1111001001100101",
    "1110101111100011",
    "0000010100011001",
    "1101110101001010",
    "1101111100100011",
    "1111101010101110",
    "1100100110101101",
    "0000010011010010",
    "1111100011010110",
    "0000010111101010",
    "0000111100000010",
    "1111101100000111",
    "0000100001000111",
    "0000000001100000",
    "0001110011100100",
    "0010000111000011",
    "1110010101011100",
    "1110100100000101",
    "1110010111011000",
    "1111110000010111",
    "1111011100011101",
    "1101110110101101",
    "0011010101010101",
    "1101100011111000",
    "0000110001001000",
    "1111111101001100",
    "1111010010001011",
    "0001101000001000",
    "1111001001000100",
    "1110111101100000",
    "0000001010000000",
    "1110110100100100",
    "0000110101101010",
    "1110010101101111",
    "0001011010111010",
    "0001100000010111",
    "0010100100111000",
    "0011000100000100",
    "0001001110010110",
    "0000111001011101",
    "1111000101010110",
    "1110011001001110",
    "1111011011101110",
    "1101101000101001",
    "1111111011110011",
    "1111000111010110",
    "1110000110111100",
    "0000111001100101",
    "1111110000100101",
    "0001101011111110",
    "0000010100110011",
    "0000001111001100",
    "0001011000110001",
    "0000010100111111",
    "1111011101010110",
    "1111001111101011",
    "1101000001110001",
    "1110110011100100",
    "1111000100110110",
    "0000000111110101",
    "0001010110010100",
    "1111001011001011",
    "0011111010001001",
    "0000001100001000",
    "0001111001000101",
    "0000001001010001",
    "1110100110100101",
    "0000111000011001",
    "1110110000010011",
    "1110010000100101",
    "1110001000111001",
    "1101111001111110",
    "1111111001001011",
    "1111111110101100",
    "0000110111011101",
    "0000111010001110",
    "1110100011110010",
    "0010000101101011",
    "1111011100010111",
    "1111100101010000",
    "0000011001101000",
    "1101010100110011",
    "0000100110110001",
    "1111000111010001",
    "0000101110001001",
    "0000000111011001",
    "0000011001001110",
    "0001011111000011",
    "1111001010111100",
    "1111101001000100",
    "0001011010001110",
    "1101111010110101",
    "0000000001001010",
    "1100111111011000",
    "1111000101010000",
    "1100011100001000",
    "1101111010101011",
    "1111111000011111",
    "1110111001111101",
    "0001000100001000",
    "0000111100111100",
    "0001110111010100",
    "0000101111001100",
    "1110110000001111",
    "1110000110100011",
    "1110111001101110",
    "1100110111000110",
    "0000001110001010",
    "1111100111100101",
    "0000110001101011",
    "0000001001001111",
    "1110011011111101",
    "0011011101011100",
    "0010000111100001",
    "0000111101110010",
    "1111011000011100",
    "1111111101101000",
    "1111100110010011",
    "1101101110101010",
    "0000010001000000",
    "1110010010010101",
    "1101000011000000",
    "0001101110101101",
    "0000010100100010",
    "0001010111110111",
    "0001110001100011",
    "0001000000001001",
    "0010010001111001",
    "1110011011110110",
    "0000011110110100",
    "1111100011010111",
    "1101101100011000",
    "1110111111110110",
    "1111011010011000",
    "0000000001001010",
    "0000111001000011",
    "1111010001100100",
    "0000011100110001",
    "0000001111010010",
    "0000110010000110",
    "0001100100100010",
    "1111100100010010",
    "0001001111101001",
    "1101011100110011",
    "1110011100010110",
    "1110011001110001",
    "1111100000000110",
    "0100000110010010",
    "0000101001011100",
    "0000100000010011",
    "0010000111010100",
    "1110110010101010",
    "1111111000100111",
    "1111101110001001",
    "1110111001001101",
    "1111101100100000",
    "1111100110110000",
    "0000100101111001",
    "1111101100011110",
    "1110110001000010",
    "0001100000011010",
    "0010001101001011",
    "0010100010101001",
    "1110100001101100",
    "0000101001000100",
    "1111110111110011",
    "1111001001011111",
    "0000100110100110",
    "1110100110101011",
    "1111000000111111",
    "1111000100101000",
    "1110011010100000",
    "0010001010011010",
    "1110000100010010",
    "0001000100100000",
    "0001100011000101",
    "1111010001000110",
    "0001110010010100",
    "1110111011101011",
    "1110101110111100",
    "1111100010100110",
    "1101111011100100",
    "1111110001111111",
    "1110000011011101",
    "0000011011101111",
    "1110111111111011",
    "1111101010110100",
    "0001011101001110",
    "1111001001111100",
    "0001011111110110",
    "1111101000110011",
    "1111010011100101",
    "0001001010101011",
    "1110000010101100",
    "1111101010000011",
    "0000010011111010",
    "1110111011000011",
    "0001110110011001",
    "1110101010000101",
    "0010011000110101",
    "0000010010011100",
    "1110000101110101",
    "0010101100011001",
    "1110111100001110",
    "0000000111101110",
    "1111000001000001",
    "1101001011011010",
    "1101000111100011",
    "1111011001000100",
    "0000000101011101",
    "0000101001011100",
    "0000011110010001",
    "0000100101001010",
    "1111010101101000",
    "0001111111100000",
    "0000111110000100",
    "1101011110111110",
    "1101111111001110",
    "1101101000001011",
    "1111100101111110",
    "0000100111010011",
    "1111000110001111",
    "0000001011111101",
    "0000001110011110",
    "0000000110101111",
    "0000010100010001",
    "1111010001000010",
    "0000000101000110",
    "1110101110111001",
    "1110110001011001",
    "1111000101111111",
    "1101101111001000",
    "1111110010000000",
    "1110010000110000",
    "0001100110101111",
    "0001011101001000",
    "0000001000000110",
    "0000100010000111",
    "1110011100010000",
    "1110111000010101",
    "0010111110100010",
    "1111101111001101",
    "0000011100101011",
    "1101001110011000",
    "1110001110111010",
    "0000001110000010",
    "0000100100011001",
    "1111100111011010",
    "1111011110000111",
    "0001001100011000",
    "1111010010010010",
    "0000110000101110",
    "0000111001001111",
    "0000111010100111",
    "1111010001111110",
    "1111110010011101",
    "1101000011100111",
    "1111100100001111",
    "1101100110001011",
    "0000110000111011",
    "0010001001011001",
    "1111011110010100",
    "0010011011111011",
    "1111100100000010",
    "0000111100100111",
    "0001100100010111",
    "1110111000101011",
    "1111001001110111",
    "1101010101111000",
    "1111001101011010",
    "1111011110101110",
    "1110001000110100",
    "0001011111010110",
    "0001001011111100",
    "0001000001101100",
    "0001000100101011",
    "1101101101111111",
    "0000100010001101",
    "1101100111000100",
    "1111010010010001",
    "1111111001111010",
    "1111101110001110",
    "0001111111010101",
    "1110101001100000",
    "0000000011010011",
    "0001101010011001",
    "0000100011101011",
    "0010110000111110",
    "0000110110000111",
    "1111010111010101",
    "0000111010011000",
    "1110101011000111",
    "1111011011100100",
    "1101100000010110",
    "0000101010010010",
    "1110110111001010",
    "1101110001000101",
    "0001100001100001",
    "0001111011100100",
    "0001010011011010",
    "0001100101100000",
    "1110111110110101",
    "0010111110111011",
    "1111001000001111",
    "0000001100111010",
    "1110011011010110",
    "1111000011011001",
    "0000100101001000",
    "1101100110111111",
    "0000011010010110",
    "0000011001001111",
    "0000001011010011",
    "0001101111111110",
    "1111111000001010",
    "1111110011111110",
    "0000000011000111",
    "1111100010000010",
    "0001111011111000",
    "1101000010011101",
    "0001110000011011",
    "0001001100101010",
    "1111001011000001",
    "0001000000100000",
    "1111001110001010",
    "0010000111000100",
    "0000100101010100",
    "1111011101010100",
    "0010001100010101",
    "1111011100001000",
    "0000100100011000",
    "1111111000100101",
    "1101110011000100",
    "1111101011010110",
    "1111100011111100",
    "1111101100110110",
    "0010000010000001",
    "0000110110111010",
    "0010010010011011",
    "0000000100100001",
    "0001001101011110",
    "0011111001100000",
    "1110101001110010",
    "1110101000100110",
    "0000000111010011",
    "1111111111010011",
    "1111000001100001",
    "0001100111101111",
    "0001110111000010",
    "0000001101101101",
    "0000011111111111",
    "0000001101100111",
    "1110001001101101",
    "0000111000101101",
    "1101111100110101",
    "0000010100011100",
    "1111000011111100",
    "1111111101111100",
    "0001101100111010",
    "1110111011011110",
    "0000000101101101",
    "0001111111110100",
    "1110111010111100",
    "0010101011000111",
    "1111011001011111",
    "0000011100011101",
    "1111101100110011",
    "1111010101110100",
    "1111011010011011",
    "1101001000101010",
    "1111111011101010",
    "1111001111111000",
    "1111010111011000",
    "0000111101010000",
    "0000001100001000",
    "1110101101101001",
    "0001101111100101",
    "0001110001100000",
    "0010010110010011",
    "1111111010100010",
    "1111011011101001",
    "1111100011110111",
    "1110011100010111",
    "0000010010011001",
    "1101111011110101",
    "0000000001010000",
    "0000101010111001",
    "1111100101100011",
    "0010110101100100",
    "0010100110110001",
    "1111100001011000",
    "0000100000000001",
    "1101010100101010",
    "0001011111100101",
    "1111100110111110",
    "1101101101111000",
    "0001100111011000",
    "1101111010110100",
    "0001100010010011",
    "0001000001001101",
    "0001011011001100",
    "0011100100101100",
    "0010101011000011",
    "0001011100101000",
    "1101000110001011",
    "1111010011101000",
    "1110100010000000",
    "1101011011110010",
    "1111000100000011",
    "1110110101111111",
    "0010011110101000",
    "0000001000010000",
    "1111110010010111",
    "0011001010101010",
    "0001010001111011",
    "0001010101001001",
    "0001011001011101",
    "1111101000101101",
    "1111110011110011",
    "1110101000001011",
    "1111000101001000",
    "1110110001011001",
    "1111101000110111",
    "0001011000000110",
    "1111101110111010",
    "0001100100011100",
    "0010010000111111",
    "0000010100000010",
    "0001100000001111",
    "1111010010001001",
    "1111101110010001",
    "1110100110101101",
    "1110111111000101",
    "0001100110011001",
    "1110001110110011",
    "0010010011001011",
    "0000101010110011",
    "1111110100101101",
    "0001000110100011",
    "1111010001100110",
    "1111111001000101",
    "0000101110011101",
    "0000010111001100",
    "0000101101111111",
    "1111000011011001",
    "0000101110001010",
    "1101001011000001",
    "1110110101100000",
    "0001101010011000",
    "0000101000110010",
    "1111111110010000",
    "0000010001011001",
    "0000101101011111",
    "0001001100010100",
    "1111100011101000",
    "1110101101100000",
    "1101101111101101",
    "1110111101011100",
    "0001011000100110",
    "0000011001011011",
    "1110110101101111",
    "1111100000100001",
    "1110100101111111",
    "0001111101010101",
    "1111011100111011",
    "0010001010001011",
    "1110111010101011",
    "1101000001011110",
    "0000011001010111",
    "1111011001000101",
    "1110100100111001",
    "1110011001111111",
    "1110110110101011",
    "1111101011000011",
    "1111111011111111",
    "0010000110110010",
    "0001011111101101",
    "1110000000101100",
    "0000110001011011",
    "1110101100111010",
    "0001011111000011",
    "0000010010110101",
    "1110001001000101",
    "0001100000000001",
    "1101101110000111",
    "0000000001100000",
    "0010010000011110",
    "0001100100011101",
    "0010101110110000",
    "0000100011101110",
    "0000010000100100",
    "0001000111011110",
    "1101111011111110",
    "0000110001000000",
    "1110011110110001",
    "0000100001001100",
    "1111001111101110",
    "1111101000111100",
    "0010000110100011",
    "1111000001011000",
    "0001011011110001",
    "0010110111111111",
    "0000000010000101",
    "0001000000000010",
    "1111011101011101",
    "1111011001011000",
    "1111110100101000",
    "1110000100000111",
    "0000001011000011",
    "1111001110011110",
    "0001101110111111",
    "0001010010111111",
    "0001101101110011",
    "1111111110001100",
    "1111100111100011",
    "0001000101001011",
    "1111100010010110",
    "1101011111010100",
    "0000110011101110",
    "1110110011111100",
    "1111101010110011",
    "0000000100010010",
    "1110001000100001",
    "0000110011111011",
    "1111110100000011",
    "0000100101110000",
    "0001100111000000",
    "0010010010010000",
    "0000110100111011",
    "1111101001101011",
    "1110101000110010",
    "0000101110000000",
    "1101001110101101",
    "0000011001100101",
    "1110001001011001",
    "0000111000100100",
    "0000110110110011",
    "0000000001011111",
    "0100111100101111",
    "1111011011111111",
    "0000110011000100",
    "0011000011100001",
    "1101100111100101",
    "0000101111100111",
    "1101000111110101",
    "0000011010001111",
    "1111111111111100",
    "1111101001111110",
    "0001000001111100",
    "0000001010100100",
    "0010110000000000",
    "1111000000001010",
    "1110010010010110",
    "0001101110010111",
    "1110010110010101",
    "1111011000000001",
    "1101111000011110",
    "1101010010110100",
    "1111110010010111",
    "1110000010100001",
    "1111100000010110",
    "0000011011000101",
    "1111000111111110",
    "0011010101111000",
    "1111000101000011",
    "0010101010011011",
    "1111111111110101",
    "1101010100000100",
    "1111100100101000",
    "1111001000100010",
    "0000011011110110",
    "1111110101001111",
    "1111010010101000",
    "0001111100010010",
    "1110011101100000",
    "0000101100100010",
    "1111011100101001",
    "1111011110001001",
    "0010010000100010",
    "1111101110001001",
    "0001111101011010",
    "1111100010111100",
    "1100000010101110",
    "0001111000010110",
    "0000000011000010",
    "1111110010100000",
    "0001000100010100",
    "0000110110001100",
    "0010011000101000",
    "0000110000111000",
    "0000101110110111",
    "0000010101010100",
    "1110110110100111",
    "1111011001101100",
    "1111100111110011",
    "1111011000101011",
    "0000010110111011",
    "1110001001100001",
    "0000001110111110",
    "1111110101000100",
    "0001000001100110",
    "0010011110001111",
    "0000100001101011",
    "0001110110011000",
    "1101100011110000",
    "1110101101000011",
    "1111100101001101",
    "1101110110011110",
    "0001011110110010",
    "0000000110110100",
    "1111110010101000",
    "0001101110000101",
    "0001011101100111",
    "0010010100100011",
    "0001101100001101",
    "0001111010000100",
    "0000100101100000",
    "1111101001000110",
    "0000011000101011",
    "1101110010001011",
    "1111101111001110",
    "1111101101010011",
    "1110101000111001",
    "0011000101001000",
    "0000001001000010",
    "0100000000100001",
    "0000111110110100",
    "0000011110111111",
    "0010111001000100",
    "0001101110111010",
    "1111111110011010",
    "1110100101101100",
    "1111000000001001",
    "1110110111110000",
    "1110011111011101",
    "0000101001001100",
    "0010010101011010",
    "0001100000010010",
    "0001111110001111",
    "0000111111011100",
    "0000100001100001",
    "0001000010000111",
    "0000101011100011",
    "0000010110010000",
    "1101111001100000",
    "1110111000010001",
    "0000011000110110",
    "0000010101110100",
    "0011011011110101",
    "1111111110010101",
    "0001011100001101",
    "0000101001010001",
    "0001100010000011",
    "0001001110111101",
    "1110100001111100",
    "0001110110110001",
    "0000001100000111",
    "1110111010100101",
    "1111001011110111",
    "1111001100110000",
    "0000111001000101",
    "1111110000001011",
    "1111110101110111",
    "0001100110000101",
    "0000100110000110",
    "1111110101101000",
    "0001011101100000",
    "0000100011001101",
    "1111111000110010",
    "1110001100001011",
    "1111111000101101",
    "0000110111111111",
    "1111100001101001",
    "0001101101001100",
    "1111011011111111",
    "0001000010111101",
    "0001111001000001",
    "0001100110100101",
    "0001111000001010",
    "1101110011000011",
    "0000000110101101",
    "1111010010011000",
    "1101111101000111",
    "1111111110001100",
    "1101111000101011",
    "0000000011010001",
    "0000000011111000",
    "1111101100111101",
    "0010000111100000",
    "0000001111011110",
    "0000101000010001",
    "0000001110000010",
    "1110110011001000",
    "0000101001100011",
    "1111011110110000",
    "1111111111111101",
    "1111011000101001",
    "1111100110100000",
    "0001000100000100",
    "1110001000111010",
    "1110111011100011",
    "1111100100000110",
    "1111101011101101",
    "0000101100001000",
    "1110010010001001",
    "1111101101100101",
    "1110101110000110",
    "1101100100011000",
    "0000110011001111",
    "1111100011000011",
    "0010110011101111",
    "0001001001011011",
    "0000001000000010",
    "0001011011010000",
    "1111110111110100",
    "0000110010110110",
    "1110100111011011",
    "1110100000100000",
    "0000111100001100",
    "1101101000001101",
    "1111110111111010",
    "0000101010011100",
    "0000000101001011",
    "0010000101100000",
    "1101101010010000",
    "0000101101101001",
    "0010001011011110",
    "0000010100001001",
    "0001010100000110",
    "1111011100001100",
    "0000110011010100",
    "1111100010000111",
    "1101011100001011",
    "0000000000101100",
    "1110100011101011",
    "0001010001001100",
    "0001010000011101",
    "0000100111010110",
    "0010001001011110",
    "1111101101001000",
    "0000111001111111",
    "0000100101101011",
    "1101010111100000",
    "0000010111101011",
    "1111001000000110",
    "1111010001001110",
    "0001001111100111",
    "1111100100000111",
    "0000111000111000",
    "1111110001000010",
    "0001000000001010",
    "0001100001001101",
    "0000101011001011",
    "0001000001000110",
    "1111011101100101",
    "0001011011010101",
    "0000010011111001",
    "1111000001100011",
    "1111011000000101",
    "1110001110110010",
    "0000100111010100",
    "0000101111101000",
    "1110011100010011",
    "0000011111000101",
    "0001000101111111",
    "0000000101100011",
    "0010011100110100",
    "1100100010110001",
    "0000101000111100",
    "1110001100110001",
    "1110100111111000",
    "0000000100110111",
    "1110001101011011",
    "0010001010110011",
    "1111111111001010",
    "1111101000110110",
    "1110110110100101",
    "1111101000101110",
    "0010011101000111",
    "1111001011110101",
    "1111101110011101",
    "0000000100010010",
    "1100110011100011",
    "0001100111011101",
    "1101110111110001",
    "0000011010001110",
    "0000011110110011",
    "0000001101111000",
    "0000000011100011",
    "0001100101110101",
    "0001011001000000",
    "0010011000011100",
    "0000001011101001",
    "0000001100111101",
    "1101010000101000",
    "1101101000111111",
    "1111101100000100",
    "1111001110010000",
    "0010010110101101",
    "1110111110000001",
    "0010000100101001",
    "0001010110010110",
    "1111001001010111",
    "0010000101010101",
    "1111010001001111",
    "1111011011111100",
    "0001010000011011",
    "1110110011101110",
    "0000000101001011",
    "1111000010101111",
    "0000011101010111",
    "0001000001001100",
    "0000100001010110",
    "0001011001011000",
    "1111010001010011",
    "0001001101001010",
    "0010010000011100",
    "1110011101010110",
    "1111001011011010",
    "1101111101011101",
    "1110111001010011",
    "1111010110000010",
    "1111011110101010",
    "0001001011011101",
    "1111010100110110",
    "0000110101010111",
    "1111111101001000",
    "1111000011111000",
    "1111111001010110",
    "1110011111001101",
    "1110100101100010",
    "1110101011000001",
    "1101111001011011",
    "1110111111011001",
    "1110101111101111",
    "0000101101100101",
    "1111111000011011",
    "0001001011100110",
    "0000011010011111",
    "1111101011001111",
    "1111010111000011",
    "0000000001101111",
    "1101011100010000",
    "1111100111011100",
    "1101011101010101",
    "1110001100011100",
    "1101100110110101",
    "1111100100011001",
    "0011010011110010",
    "0010001001001011",
    "0000110010010001",
    "0001001110110101",
    "1111011101000100",
    "0001011000101001",
    "1110000101011011",
    "1101110000001001",
    "1111010101111100",
    "1100111110010100",
    "1110010010011110",
    "0001001000111011",
    "0000001000110111",
    "0001001111111011",
    "0001010000101000",
    "0000010100001011",
    "0000011110110000",
    "0001010110001100",
    "0000011101000111",
    "1110111011000101",
    "1111101010011100",
    "1110111011000000",
    "1110100001111000",
    "1110111000000001",
    "1111101110101010",
    "0010111111101110",
    "1111100010001001",
    "0000110001011100",
    "0001101011111001",
    "0000111111100000",
    "0010010001101111",
    "1111010001100001",
    "1111000010011000",
    "0000000000100101",
    "1110000111101010",
    "0001100100010110",
    "1101010110110110",
    "0000100000110101",
    "0010001000100111",
    "1111100100101000",
    "0001011000000001",
    "1111001000100011",
    "0000100100001111",
    "0000001010111110",
    "1110111001101110",
    "1111010011101100",
    "1110010010000001",
    "1110110001101000",
    "1111010011011001",
    "1110001010100110",
    "0001000001101101",
    "0011011111010110",
    "0100101011110110",
    "0010011011001011",
    "0000101101010001",
    "0000000001111110",
    "1110011010110100",
    "1111000011010110",
    "1111111010100010",
    "1110101011101001",
    "0000010011001011",
    "1110011011001100",
    "1111011100100011",
    "0000110110011010",
    "0001001101001110",
    "0010011011010110",
    "0000001111111001",
    "0001100000001010",
    "0000111101001100",
    "1101001001100001",
    "0000001101011011",
    "1101110001011110",
    "1101010110000110",
    "1110010101111101",
    "1110101011110001",
    "0010001000100111",
    "1111101100001101",
    "0001100010100011",
    "0000011000010011",
    "1101110000110100",
    "0001011001110010",
    "1110000011010111",
    "0000110110000010",
    "0001000111010100",
    "1101110100111100",
    "0001011000100100",
    "1111101110000000",
    "1110111101001111",
    "0000110011111100",
    "0000010101000001",
    "0010100001011110",
    "0000101111101000",
    "0001100001001111",
    "0001000011001110",
    "1110011100111110",
    "0000100100100000",
    "1011111100100011",
    "1110001101100000",
    "0000110111111010",
    "1110010101111100",
    "0001101000101111",
    "0001011011011001",
    "0000011000111000",
    "0000010100011000",
    "1111011011010110",
    "0001110000000000",
    "1110110011001000",
    "1110101100011010",
    "1101110011100111",
    "1101110101000010",
    "1111111110000100",
    "1110001110101110",
    "0000000111000010",
    "1111101111111110",
    "0000100111011101",
    "1111110100110101",
    "0000001101100100",
    "0001100000111001",
    "1111100001011110",
    "1110101101010100",
    "0000011110111001",
    "1101100101011001",
    "1111010111011001",
    "0000000101010111",
    "1110000100010000",
    "0010001001001111",
    "0001000000111011",
    "0001100110010101",
    "0001010010101111",
    "1110110000010110",
    "0001110011011101",
    "1101110010011011",
    "0001010000110011",
    "1111111001111110",
    "1110011101101011",
    "1111110011000010",
    "1100100101101100",
    "1111001011010010",
    "0001001101011101",
    "0010011110101101",
    "0010101111011000",
    "0000011000001000",
    "0000010011011001",
    "0000011111101000",
    "1111101110100100",
    "1111111011111110",
    "0000000101110011",
    "1110001010001011",
    "1111010010111010",
    "1111000011100110",
    "1111010110101110",
    "0000011111000100",
    "0001010110110000",
    "0001010110111100",
    "0000101101101111",
    "0010010110100101",
    "1111110011100101",
    "1111001100111111",
    "1111010101010011",
    "1110100011010110",
    "1110111011110010",
    "1101101110101011",
    "1111111100011110",
    "0000111011000011",
    "0001110110111011",
    "0010110011000010",
    "1111100111111111",
    "0000001101110100",
    "0001111001111101",
    "0001011111111011",
    "0000010110111100",
    "1101101110000101",
    "1101111101110111",
    "0000101001011000",
    "1111010010110001",
    "0010011110010111",
    "1111000000101110",
    "0001100001001010",
    "0000100111111010",
    "0001001100011110",
    "0000110000100000",
    "1110111010101001",
    "1111010100101110",
    "0000010111111001",
    "1110101000001001",
    "1111001011111101",
    "1110001000011111",
    "1111010100111000",
    "0001010110011100",
    "0000011001100011",
    "0000010111010101",
    "1110001010010001",
    "0000110011011111",
    "0001000100011011",
    "1110111011110010",
    "1110101001011011",
    "1100101001011010",
    "0000001111110001",
    "1111100001101011",
    "1110100111100001",
    "0010101000000001",
    "1111000111111010",
    "0001011010011100",
    "0001101100100000",
    "0000101111010110",
    "0000011101000110",
    "1111010111000110",
    "0010011010111001",
    "1101110111011100",
    "1110101000100000",
    "1111111101100001",
    "1101111100000011",
    "1111100010100011",
    "0001010101111100",
    "0010011000100000",
    "0001001101001100",
    "0000100110111011",
    "0000010010010011",
    "0010010110010011",
    "1111010011110101",
    "0000000011011001",
    "1110110100011010",
    "1111010111111011",
    "0000110001110110",
    "1110110100010111",
    "0000001100000000",
    "0000001010101010",
    "0010110101101011",
    "0000000101001100",
    "1111101011010111",
    "0010010100000110",
    "1101000101010110",
    "0000010011000001",
    "0000001000011101",
    "1110011010011001",
    "1111011010111011",
    "1110110000100001",
    "0000011101110001",
    "0001110001111011",
    "0000101110110001",
    "0001101001100101",
    "0001101011111111",
    "0000110010110100",
    "1111100011110010",
    "1110010100111011",
    "0001000011001011",
    "1110011001001110",
    "0000010001001010",
    "1111101111011010",
    "0001011111011001",
    "1111101001001011",
    "1111100000010000",
    "0001001100011000",
    "0001010111011111",
    "0001011000000101",
    "0001100001110101",
    "1110111000111000",
    "1111101111011000",
    "0000001000010111",
    "1101100000100111",
    "0000101001000101",
    "1101001100110100",
    "0000010010110000",
    "1111111001110011",
    "1111011010100001",
    "0010010010000101",
    "1110111100010011",
    "1111110110110010",
    "1110110110110010",
    "1100100010010110",
    "0000000010100010",
    "1111010111001001",
    "1111001100101000",
    "1111011100000001",
    "1101111101001111",
    "0010111001000111",
    "1111101010111011",
    "0010100100100101",
    "0001101000111100",
    "1111101010000011",
    "0010011001000010",
    "1111111111000111",
    "1111100011110110",
    "0000101011001110",
    "1111111110101111",
    "0000001000000010",
    "1110100000100111",
    "0000110001101100",
    "0001001100100101",
    "0000110111111111",
    "0001101111101001",
    "0000110010000101",
    "0001111001001100",
    "0000100011001010",
    "1110111010110010",
    "1110111011111101",
    "1101000001101011",
    "1101111010101111",
    "1110011011010110",
    "1110110110010011",
    "1111101100011011",
    "0010001010101000",
    "0010000001000101",
    "1111001101011100",
    "1110110000111111",
    "0001001100111011",
    "1101010010100111",
    "1111001101100011",
    "0000011110000110",
    "1110000010001111",
    "0000000111111011",
    "1101110000111000",
    "1111110100001111",
    "1111011111100101",
    "0000011011100111",
    "0001100011000100",
    "0000110110011100",
    "0010000101010000",
    "0001011100101111",
    "1110101110110000",
    "1111101011111110",
    "1100111110011001",
    "1111011111110111",
    "0000101000011001",
    "1110101010011010",
    "0001001000101100",
    "0000100010010100",
    "0010001001000100",
    "1111110111000101",
    "0000000111101011",
    "0001100000010100",
    "1110110110100100",
    "0000100100001000",
    "1111000000111110",
    "1101010111110110",
    "0000011101111001",
    "1111001110011010",
    "0000001001111000",
    "0001101001000001",
    "1110100011001010",
    "0000111011001101",
    "1100111111101100",
    "0001010111011100",
    "1111011000011000",
    "1110100000110001",
    "0001001100110100",
    "1110010000000000",
    "1110111100000101",
    "1110110100101100",
    "1110110000110110",
    "0001111010010111",
    "1110011001110110",
    "0001001101011001",
    "0010000011110110",
    "1110011111111101",
    "0001111110100111",
    "1111101011111101",
    "1110110010100010",
    "1101110111111111",
    "1110101000011101",
    "0000111111111101",
    "1111010110000010",
    "0001001000101000",
    "1111101010011010",
    "0000101001101011",
    "0001011010111000",
    "1111100000011000",
    "1111010010100000",
    "0001011110001101",
    "1110111100001011",
    "0001001100011101",
    "1111101101011100",
    "1110001111011111",
    "0000010100001001",
    "1110111111011010",
    "0010001110010011",
    "0001000001110001",
    "0010000110010010",
    "0000011101011100",
    "1111110010110010",
    "0001100100101100",
    "0010001010011000",
    "0000111001011111",
    "0001101100110011",
    "1110100111010000",
    "0000011001110010",
    "1111011000001110",
    "1111110110000001",
    "0010000101100010",
    "1111111010001110",
    "0000101000000110",
    "0000111100000011",
    "1111010001101100",
    "1110100001110001",
    "1111000011011100",
    "1111001111010111",
    "1101010010011100",
    "1111001101111010",
    "1111001011101100",
    "1110110001111110",
    "0001100101001100",
    "1110110000000110",
    "0000000011011011",
    "1111001011011010",
    "1111100001111010",
    "0001111110010011",
    "1110010011010010",
    "0000001011000100",
    "1111111010110110",
    "1111001100001001",
    "0001001011100011",
    "1110000100111001",
    "1111100000111101",
    "0000111001001011",
    "1111011001110000",
    "0011011100111110",
    "0001011100100111",
    "0000111100001010",
    "1111111100011101",
    "1111010001101011",
    "1111100010001110",
    "1110000100101110",
    "1110110110010101",
    "1111110001101111",
    "0000001000011100",
    "0010000011010011",
    "0001000100000100",
    "0000010111001110",
    "0001011101010010",
    "1110111011111100",
    "0001101100011010",
    "1111010101000101",
    "0000111101111101",
    "0000011110101000",
    "1110110110100010",
    "1111101011111001",
    "1110010010100001",
    "1110010100100000",
    "0000011001011000",
    "1110100001000010",
    "0010111011100001",
    "0000111110000010",
    "0000111110111011",
    "1111111111100101",
    "1110111010001000",
    "0001110010111101",
    "1111100011000101",
    "1110111011100101",
    "1111110101110001",
    "1101111000100001",
    "0001101101011011",
    "0000101010001011",
    "0010001011011000",
    "1111101111110001",
    "0000011011001011",
    "0000011100011110",
    "1110101000001000",
    "0000011101011011",
    "1111101011010111",
    "1110000010010000",
    "0000110011000011",
    "0000011001100101",
    "1111101111111001",
    "1111011111101010",
    "1110111001111011",
    "0001000011100100",
    "1111011001010110",
    "0001011010111111",
    "1110010010010100",
    "1111000000000101",
    "1111011010011010",
    "1111010011000110",
    "1110100001100001",
    "1111101011011110",
    "1110000100001110",
    "0000101000001010",
    "1111101010001111",
    "0001000011001000",
    "0000110000001011",
    "0001000011000110",
    "0001110110111111",
    "0000110110111101",
    "1111011001001111",
    "0000011100100010",
    "1100000110011000",
    "0000110101000101",
    "1111001000110000",
    "1111111111110110",
    "0001100010100101",
    "0000111100011110",
    "0011000010001010",
    "0000011111001011",
    "0001011100100010",
    "1111101100101010",
    "1101101010111000",
    "1111111011000110",
    "1110011000101011",
    "0000010101001000",
    "1110111000011001",
    "1110100000111010",
    "0100010010001001",
    "1111010011000010",
    "0011001100101011",
    "0010001111010010",
    "1111010111001011",
    "0001001100111101",
    "1110110010011101",
    "0000001001010010",
    "0000101111101011",
    "1100100011111010",
    "0010001101101111",
    "1111100010110000",
    "1111110100101011",
    "0000101110000000",
    "0000010111011111",
    "0010010010111101",
    "0001010001001010",
    "0001111011110110",
    "0000000000110110",
    "1110101000101010",
    "0000111011001100",
    "1110010100011011",
    "0000100001000000",
    "1110111111000010",
    "1111011110011011",
    "0001100110001111",
    "0001010011111101",
    "1111111011101010",
    "0001010001110100",
    "1111111110010011",
    "1110111101111001",
    "0000010000000111",
    "0010011110110001",
    "1111001001011010",
    "1110011111000110",
    "1111101110011111",
    "1111001001100100",
    "1111111111011111",
    "0000101111100100",
    "0001101011111000",
    "0001001001110010",
    "1111011111011101",
    "0000110001001110",
    "0000001111010100",
    "0000001101000110",
    "0010001110001110",
    "1101001110001000",
    "1110101111010000",
    "0000001100010011",
    "1110100111110111",
    "0011010011010100",
    "0001100011100101",
    "0001110101100011",
    "0001110101110110",
    "1111100101001110",
    "0010000100101010",
    "0000001000011001",
    "1111110100000011",
    "0001010011101011",
    "1110110111101001",
    "0000000101001011",
    "1111001000101110",
    "0001011101111111",
    "0000011100100110",
    "1111111110110110",
    "0100010111111001",
    "1111100101111110",
    "0001110010101001",
    "0001001100001010",
    "0000010110101011",
    "0000101101111001",
    "1011101110111101",
    "1110100001101101",
    "0000001011101111",
    "1111010000101111",
    "0011010001011000",
    "0001010100111000",
    "0001110001100100",
    "0001010111000100",
    "1110010111110010",
    "0011001011000001",
    "1111001000110100",
    "1110001000000010",
    "1111110100000000",
    "1110010011010100",
    "1111100111101110",
    "1111010000100010",
    "1111101010100001",
    "1111011111110011",
    "1110010100000010",
    "0001101000101110",
    "1111011100001011",
    "0001010010001111",
    "1110110111101000",
    "1110100011101001",
    "1110101011111001",
    "0000000000100011",
    "1111010000110010",
    "0000111001011101",
    "1111011111111010",
    "0010001101111011",
    "1110110001000000",
    "0010100010010000",
    "0010101110101111",
    "1101110101111110",
    "0001001000011111",
    "1110010110100000",
    "1111110101000000",
    "1110100001110111",
    "1110011110100110",
    "0000110010011100",
    "1111000000101001",
    "0000010000001110",
    "1111100011100011",
    "0000000111111111",
    "0001011110101010",
    "1110110010011101",
    "0000110010011110",
    "0000001010011000",
    "1110111101010001",
    "0001001011101111",
    "1110110001100111",
    "0000101011110110",
    "1110111100010100",
    "1110001000111001",
    "0001001101101101",
    "0001010011011010",
    "0010100101001101",
    "0001001001101110",
    "1111010100101011",
    "1111110010011101",
    "1111101011001111",
    "1111101100011100",
    "1110001100111001",
    "1101110111010100",
    "1110010111001001",
    "1111001100100000",
    "0000001100101010",
    "0010011110011110",
    "1110101101010011",
    "0010111110000111",
    "0000001101100000",
    "0000111011010111",
    "0001000101101010",
    "1111111101010111",
    "1111000111101011",
    "1111100001001001",
    "1110001010110101",
    "1110100110001111",
    "1110010101001100",
    "0010000010111010",
    "1110110110011010",
    "0001100111001100",
    "0001101100001000",
    "0000000100101111",
    "0001110111010001",
    "1101110101001011",
    "0000101011011110",
    "1111011111100010",
    "1110111011011101",
    "1111001101010010",
    "1110110100010011",
    "0001001111111110",
    "0001110110111110",
    "1111111110111010",
    "0000001001011000",
    "1110111110000111",
    "0001000100000100",
    "0001001010101000",
    "1111001110100111",
    "1111100101000001",
    "0000011100011000",
    "1111011100111010",
    "0000100010011000",
    "1110100101101000",
    "0000001100011011",
    "0000100110101111",
    "0010010100001011",
    "0011000110011001",
    "1111011001000001",
    "1111101011100110",
    "0000100111101111",
    "1111111011111001",
    "1110010000001001",
    "1101101000111100",
    "1111011000011101",
    "1111111011010010",
    "0000111101101100",
    "0001000101100111",
    "0000010011101101",
    "0001001011011011",
    "0001000011110111",
    "0001001100001111",
    "0000000111000101",
    "1110100101001010",
    "0000000101101110",
    "1101010011111101",
    "0000000111101110",
    "0001000100000101",
    "0001011110100100",
    "0001110100000010",
    "1111000110001111",
    "0001011110101000",
    "0000010001010100",
    "1111010011101001",
    "0000101001100111",
    "1110001010111010",
    "0000000011001100",
    "1110010000111001",
    "1110110111011100",
    "0000111111001000",
    "1111110011011000",
    "0000010110011111",
    "0001011101101100",
    "0001110111101101",
    "0010000011011001",
    "1111111000111011",
    "0010100111100001",
    "1101110111001111",
    "1110010011110000",
    "0010100111110001",
    "1101101110100011",
    "1110110100011010",
    "1110011100011111",
    "1111110010111111",
    "1111001100101111",
    "1111000111101110",
    "0001110110000011",
    "0001010001101011",
    "0000100010110100",
    "0001011011111000",
    "1111101011110100",
    "1110011000100110",
    "1111100110001111",
    "1100101000011110",
    "0000111110010111",
    "1110011101000110",
    "0001000001101111",
    "0000010011101011",
    "0000011001010110",
    "0011000011011101",
    "1110000101100111",
    "1110111110100100",
    "1110100010100010",
    "1111100111010010",
    "0000100110001010",
    "1101011111110001",
    "0000111000001101",
    "1111110011110011",
    "1101011010101011",
    "0000010010100011",
    "1110100010001110",
    "0010001110111000",
    "0000101011010011",
    "1110101111111000",
    "0000101110110110",
    "1110001010101101",
    "0000100001100101",
    "1111110110110101",
    "1110100000000101",
    "0000100110110101",
    "1110110011101110",
    "1111011011000100",
    "0001011000101111",
    "1111001111110000",
    "0000111011011001",
    "1110111111100100",
    "0001101101101110",
    "0001010110100101",
    "1101000000011010",
    "0000000010110000",
    "1110011100110111",
    "1110110001001101",
    "0000011011101100",
    "1111010000100001",
    "0001001010000000",
    "1111010111001101",
    "0001111101000110",
    "0010001000001000",
    "0000011000111010",
    "0001000100011100",
    "1111111011001011",
    "1110110000111100",
    "1111100001100001",
    "1111100110000110",
    "0000000000000101",
    "1101111010111110",
    "0010010100001011",
    "0000100110010001",
    "0000100000100100",
    "0001001100100100",
    "0000010110101110",
    "0001010011111101",
    "0000011000000110",
    "1111000101110110",
    "0001011001010100",
    "1100110010110111",
    "1111100101011011",
    "1101101011100011",
    "1111000010000011",
    "0011001111010101",
    "0000110111000111",
    "0001010001010101",
    "0000111100001000",
    "0000011100101100",
    "0010010111011011",
    "1111000001001011",
    "0001010010010101",
    "1110100100000100",
    "1100001100111000",
    "1111011100010110",
    "1110100100001110",
    "1111111111111100",
    "1111111111110110",
    "0001011001111001",
    "0000011000100100",
    "1111100100110101",
    "1111111000000010",
    "1111111001011101",
    "1110000110010110",
    "0000101010110110",
    "1101001010000110",
    "1110100011110000",
    "1111110001011101",
    "0000000101100111",
    "1111011101000110",
    "0001101110000100",
    "0000011001100011",
    "0001111011001110",
    "0000111110000011",
    "0010101000011101",
    "1110011111001000",
    "1111101100100010",
    "1111001101111000",
    "1101100101111110",
    "0000011101100111",
    "1111000111111011",
    "0000000001010000",
    "0000111110100011",
    "0010101111011011",
    "0001111111100001",
    "0000110001110001",
    "0000011000011110",
    "1111110110000001",
    "1110011010110110",
    "0000110000010111",
    "1101011001011011",
    "1101100001101100",
    "1111101110011001",
    "1110100100010011",
    "0001100101101101",
    "0000000000010011",
    "0010000000011100",
    "0010001011011011",
    "1110100110000010",
    "1111110010001101",
    "1111100000011001",
    "1111111110100110",
    "1110011100001011",
    "1111011011111011",
    "0000001110010101",
    "1110111000111000",
    "0000101001010101",
    "0001100110010110",
    "0001100101111000",
    "0001101111001111",
    "1110010101100011",
    "0001110110111100",
    "1111011100011011",
    "0000000000100100",
    "1111100110100000",
    "1111101100001100",
    "1110100100101100",
    "1110100011110010",
    "1111111101011110",
    "1111111100100011",
    "0000100110011100",
    "0001101101110010",
    "0001001000100110",
    "1111100101000001",
    "0011010111011111",
    "1110101000010001",
    "1111011110110100",
    "1110011100001100",
    "1101011000101011",
    "1111100110111000",
    "0000011110011000",
    "1111111110110100",
    "0000001001111010",
    "1111100111101000",
    "0010101101101110",
    "1110110000000110",
    "0001011110001101",
    "1111000010100110",
    "1110101000100110",
    "1110010111010011",
    "1110101111000010",
    "0000000100100111",
    "1110111110111111",
    "1111010100100100",
    "0001011110001101",
    "0001000101000100",
    "0001011001111111",
    "0010010100010011",
    "1111110011011010",
    "0000101010010010",
    "1110111101110011",
    "1111011110001110",
    "0000010000101101",
    "1110001001001001",
    "1111010110011001",
    "1110100111000100",
    "0001100011110111",
    "0000011011100001",
    "1111011010001010",
    "0010111110111110",
    "0000001010110010",
    "0000011110110111",
    "1111101000100001",
    "1101010010010001",
    "0000010110000010",
    "1101111000011100",
    "1111101100101100",
    "1110001101110001",
    "0000010100110101",
    "0001110010111101",
    "1110010110100111",
    "0010010101011011",
    "0000101100001010",
    "0000001110001110",
    "0001100001110101",
    "1110001000000010",
    "1100110011110111",
    "1111111010100011",
    "1101110110110110",
    "1111100101111101",
    "1111001011110010",
    "1111101011101010",
    "0001100001000010",
    "0000001101111110",
    "0001000000100100",
    "0000111001110111",
    "0001010100011100",
    "0001100111111100",
    "1101110111110110",
    "1111010010111011",
    "1110100000110010",
    "0000000010111110",
    "0000011111111111",
    "1111000000101001",
    "0001000100101100",
    "0000100100101010",
    "0011001111100000",
    "0010001010011000",
    "0000000000010010",
    "0000101111000001",
    "1111100000001110",
    "1111001100000000",
    "1111100111100010",
    "1110111110100010",
    "0001000111011000",
    "1111010110100111",
    "0001101111111111",
    "0010101100100011",
    "1110001010110111",
    "0000001110001011",
    "1111001001010000",
    "1110110110001101",
    "0000000000111100",
    "1110011011011100",
    "0000011100010000",
    "1110011111000011",
    "1110101100010111",
    "1110110110111100",
    "1111110011000001",
    "0000111011010101",
    "1110100011001000",
    "0001010010011011",
    "0001011110110101",
    "1111100000100101",
    "0001111110010000",
    "1111001110101100",
    "1111011101010111",
    "1111010101011101",
    "1110101010000011",
    "1111101111111110",
    "1101101101011101",
    "0000001101110110",
    "0000111110010101",
    "0000100100111010",
    "0001111110000101",
    "1111100111000010",
    "0001011100001111",
    "0000010000100010",
    "1111100100101000",
    "0000000110011110",
    "1110001100010101",
    "1111010010011001",
    "1110110000000001",
    "1110000100111010",
    "0000010110010001",
    "0001101101000111",
    "0001000100111101",
    "0010001101111101",
    "0000010001001110",
    "0011001010110001",
    "1111111011100100",
    "1110011100011101",
    "1111000011010101",
    "1111000101110011",
    "0000011110101011",
    "0001000001111101",
    "0000010100101111",
    "1111010010110000",
    "0000100000101111",
    "0001000101101001"
  );

  constant PKG_INPUTSAMPLESFI_CONCAT : std_logic_vector(40015 downto 0) := (
    "0010100010011010" & 
    "0001111001101011" & 
    "1110100101100000" & 
    "0001001110111110" & 
    "1111000101011000" & 
    "1110111000100010" & 
    "1101110000111111" & 
    "1111101110001101" & 
    "0011010000000000" & 
    "0001110001011110" & 
    "1111111101011001" & 
    "0010111101000111" & 
    "0010000000001100" & 
    "0001001101101111" & 
    "0000101000101000" & 
    "0001000110101010" & 
    "1110111000010010" & 
    "0001001010010101" & 
    "0000110010011101" & 
    "1111100111011011" & 
    "0000110111001101" & 
    "1101100011101100" & 
    "0001000101101101" & 
    "0010011110011010" & 
    "0000100011100110" & 
    "0011000010001110" & 
    "0000110010110101" & 
    "0000100010101010" & 
    "0000101010100111" & 
    "1101111110100110" & 
    "0001000101000101" & 
    "1101000011010100" & 
    "1110010011110111" & 
    "1110110111001011" & 
    "1100000011110011" & 
    "0010101111110101" & 
    "0000001111101100" & 
    "0000100001011101" & 
    "0010101001011110" & 
    "1110001101010110" & 
    "0001001101001111" & 
    "1110110000110010" & 
    "1111111111011010" & 
    "1111101100010011" & 
    "1101010101011000" & 
    "0000001010010011" & 
    "1110100110011011" & 
    "0000111111111110" & 
    "0001111100000010" & 
    "0001001011010011" & 
    "0001001000101110" & 
    "0000001001010000" & 
    "1111101000010111" & 
    "1111010000100010" & 
    "1110110000100010" & 
    "0001101110010100" & 
    "1101011011011110" & 
    "1111110000000011" & 
    "1111011100100011" & 
    "0000000111101111" & 
    "0000001110000101" & 
    "1111111100111101" & 
    "0001110101001000" & 
    "0010011000001101" & 
    "0001011101101101" & 
    "0001011001010010" & 
    "1101100000110001" & 
    "1110111011011110" & 
    "1110010100010101" & 
    "0000100011001010" & 
    "1111100100110101" & 
    "1111100000110110" & 
    "0000001011011111" & 
    "0001101110111100" & 
    "1111010011010111" & 
    "0000100110010000" & 
    "1110101001010010" & 
    "0001010101010100" & 
    "0000001100011100" & 
    "1110100100011011" & 
    "0001100111000100" & 
    "1110011111011001" & 
    "1111100100111100" & 
    "0001010000100110" & 
    "1110001100110000" & 
    "0010000000010111" & 
    "0000110000010101" & 
    "0001000010001011" & 
    "0001011111100100" & 
    "1110110000010001" & 
    "0000001010010100" & 
    "1111000110111100" & 
    "0000011001001101" & 
    "0001111101110000" & 
    "1101100010000011" & 
    "0000011000001110" & 
    "1110101011101100" & 
    "1110011100000101" & 
    "0000011001111110" & 
    "1110010001011101" & 
    "0010110101110010" & 
    "1111001011011110" & 
    "0000111100011110" & 
    "1111110100111101" & 
    "1111000100011001" & 
    "1111100101110011" & 
    "1110101100000101" & 
    "0000000111100110" & 
    "0001011000100011" & 
    "1110110011110100" & 
    "1111001010111011" & 
    "1111000101001001" & 
    "0010101000011101" & 
    "0000001101001010" & 
    "0000111000011000" & 
    "0001011011101110" & 
    "0000011100001011" & 
    "1101101101011111" & 
    "1111001011101000" & 
    "1100111111011011" & 
    "0011000110010101" & 
    "1111100101110010" & 
    "0001110000000011" & 
    "1111110010010110" & 
    "1111100110010100" & 
    "0001101110100100" & 
    "0001001010100111" & 
    "0000100100010010" & 
    "0001000100101100" & 
    "1100101101101010" & 
    "1111110101100101" & 
    "1101011000000001" & 
    "1101110011010110" & 
    "0000001011100000" & 
    "1111010010010010" & 
    "0001010101111011" & 
    "1110100101100001" & 
    "0010011001111011" & 
    "0001101000001011" & 
    "1111100111101111" & 
    "0001010101001111" & 
    "1110101111011110" & 
    "1101111010111110" & 
    "1111000101111111" & 
    "1101010111100001" & 
    "1111001101100011" & 
    "1101100110111110" & 
    "1111110101101001" & 
    "1110110101111010" & 
    "0001000010000001" & 
    "0010100001010010" & 
    "0000000011000010" & 
    "0000110011110110" & 
    "1111100100101110" & 
    "1111110010001011" & 
    "0000000011101101" & 
    "1101011111000000" & 
    "0000101110110001" & 
    "1111011100100110" & 
    "1110011010100010" & 
    "0001000000111111" & 
    "1111000100100111" & 
    "0000001010000101" & 
    "0011110011011100" & 
    "0001100100110101" & 
    "0001100111011101" & 
    "1101101111110010" & 
    "1110110011100110" & 
    "1111001100111110" & 
    "1110111111011000" & 
    "1110110110111110" & 
    "1100011011110111" & 
    "1110111011000011" & 
    "0001001011011011" & 
    "0000011101010111" & 
    "0010011100111010" & 
    "1111111011111110" & 
    "0001000001110101" & 
    "1111111001010101" & 
    "1111101000001001" & 
    "1110110101000101" & 
    "1110101001110110" & 
    "1110100001111101" & 
    "1111010101100011" & 
    "1111100011100111" & 
    "0010010110010010" & 
    "1110110011010110" & 
    "0010100010011101" & 
    "0001111100000001" & 
    "1111110110100010" & 
    "0001000111010010" & 
    "1110110010010011" & 
    "1111010111100101" & 
    "1111011001110000" & 
    "1110010000000001" & 
    "0001000001000110" & 
    "0000010010101101" & 
    "0000110101101011" & 
    "0000101000101001" & 
    "0000101100010100" & 
    "0010001011101110" & 
    "1111000010011010" & 
    "0001110010110100" & 
    "0000101011011101" & 
    "1110111001101000" & 
    "0000101101001101" & 
    "1110011101011101" & 
    "1110011100000001" & 
    "1111100000100110" & 
    "1110110110111001" & 
    "0000110001101111" & 
    "0001100110100010" & 
    "0000011001101110" & 
    "0000110010110011" & 
    "1111001101010100" & 
    "0000001000101000" & 
    "1110110011111011" & 
    "1111011001011100" & 
    "0000111010001101" & 
    "1101111100110011" & 
    "1111001000000111" & 
    "0000010111100110" & 
    "0001100110110100" & 
    "0000100111011000" & 
    "1110100011111010" & 
    "0001100011100011" & 
    "1111111010010101" & 
    "0001000111101111" & 
    "0000000111000101" & 
    "1111001101010111" & 
    "0000100101010011" & 
    "1100111100101100" & 
    "1110011011100111" & 
    "1110111011100011" & 
    "1110011111101111" & 
    "0000111111010001" & 
    "1111111011101011" & 
    "1110001111111010" & 
    "0000110100100001" & 
    "0001001010011001" & 
    "0000001111100001" & 
    "1111111011111111" & 
    "0000000001011010" & 
    "1111010110011011" & 
    "1110011000011010" & 
    "1110101000000100" & 
    "1110101011100100" & 
    "0001111110011101" & 
    "0000111100010111" & 
    "0000000110111101" & 
    "0001010001000001" & 
    "0000000010010101" & 
    "0001000100111100" & 
    "0000110011000101" & 
    "1110011001000111" & 
    "1111111101000110" & 
    "0000001110010000" & 
    "1101000111101111" & 
    "0001111001101011" & 
    "1111010101110101" & 
    "0010010011110010" & 
    "1110010000011000" & 
    "0000101100000000" & 
    "0000111111111110" & 
    "0000010101111100" & 
    "1111101000111001" & 
    "1111011110011011" & 
    "1110011101010111" & 
    "1111011100100000" & 
    "1110110110011111" & 
    "0000100001001010" & 
    "1111110110010001" & 
    "0001011000001100" & 
    "0000001100011010" & 
    "0000010100110001" & 
    "0001000011100100" & 
    "1110101111101110" & 
    "0001110001010001" & 
    "0000010111110011" & 
    "1110101101011101" & 
    "0001000110100010" & 
    "1110110010110010" & 
    "1111101110101100" & 
    "0000111011000000" & 
    "1111111011101111" & 
    "0001100011001000" & 
    "1111001110101100" & 
    "0000101000000100" & 
    "0010011110000100" & 
    "1110010011101110" & 
    "0001010010001110" & 
    "1101000011100000" & 
    "0000101100010011" & 
    "0000001111011011" & 
    "1110001100110011" & 
    "0000000111101100" & 
    "1100010001110110" & 
    "0000111100111111" & 
    "1110101001110000" & 
    "1101101111111000" & 
    "0010000101000111" & 
    "1111000111100111" & 
    "0001010000011010" & 
    "0001000011001000" & 
    "1111100111111000" & 
    "1111011111111111" & 
    "1110101001011111" & 
    "1111011110101110" & 
    "0000011111110110" & 
    "1111100010100011" & 
    "0010001101001111" & 
    "1111110010011100" & 
    "0001001000010110" & 
    "0010010010010001" & 
    "1101110010111110" & 
    "0000110011011111" & 
    "1101101110111010" & 
    "1111010010100000" & 
    "0000000001110010" & 
    "1111000001100101" & 
    "1111001011010001" & 
    "1110010010110101" & 
    "0000100000100100" & 
    "0000100011011001" & 
    "0000010111101000" & 
    "0010011001100110" & 
    "1111001000110010" & 
    "0000101010110000" & 
    "1110001111010110" & 
    "1111111010010010" & 
    "1111100011111110" & 
    "1100111111101100" & 
    "1111001000000001" & 
    "1110001111100011" & 
    "1110111110111001" & 
    "0000101111111001" & 
    "0010000110010000" & 
    "0010011010101000" & 
    "1110110001111110" & 
    "0000010111001000" & 
    "1111111010010011" & 
    "1110101111111010" & 
    "1111110101100000" & 
    "0000001000001000" & 
    "1101111011010000" & 
    "0001110001000111" & 
    "1110010010001100" & 
    "0000101100110000" & 
    "0001100000100111" & 
    "0000001001110001" & 
    "0010111000011000" & 
    "0000011000111111" & 
    "0000000011111001" & 
    "1110100100010000" & 
    "0000100111111011" & 
    "1111100101100010" & 
    "1110010011010110" & 
    "1111111100010100" & 
    "1111110010010000" & 
    "1110000110010101" & 
    "0000110101110110" & 
    "1111110010111001" & 
    "0010110000011011" & 
    "0000011010101011" & 
    "0000101101000110" & 
    "0001100111100010" & 
    "1110110001010001" & 
    "1110100111010101" & 
    "1111000110000110" & 
    "1110000111001011" & 
    "1110101110001100" & 
    "1110111101010001" & 
    "1111100011001011" & 
    "0000110000000010" & 
    "0000011001110101" & 
    "0001000110000111" & 
    "1111110001110111" & 
    "0001001100011110" & 
    "1110100010010011" & 
    "1111110011010010" & 
    "0010100111011001" & 
    "1111001010001000" & 
    "1111000100000100" & 
    "0000000110011010" & 
    "1101111101111011" & 
    "0011001011111101" & 
    "0000110111000101" & 
    "0010000100001010" & 
    "0000011001101101" & 
    "0000001111010111" & 
    "0000110000000011" & 
    "1110101100010011" & 
    "1111000110100000" & 
    "1110010110101000" & 
    "1101010010100100" & 
    "1111111110110011" & 
    "1101000100010000" & 
    "0000111110101100" & 
    "0000101110100010" & 
    "0000110001000011" & 
    "0010010001010000" & 
    "0000100011111100" & 
    "1111010111001010" & 
    "1111010110100000" & 
    "1110010100010111" & 
    "0000010011001111" & 
    "1111010100111110" & 
    "1111000101101110" & 
    "0000111011101110" & 
    "1111011110101010" & 
    "0010011110111011" & 
    "0000000011000000" & 
    "0000100111101111" & 
    "1111110010111101" & 
    "0000000100110101" & 
    "0010001000001011" & 
    "1110101101100000" & 
    "1111001000011000" & 
    "1111000100100001" & 
    "1101000110100011" & 
    "1111101100101011" & 
    "1110100101011010" & 
    "0000011010101111" & 
    "0000110001111111" & 
    "0000101011011100" & 
    "0010000111000000" & 
    "0001111000011010" & 
    "0001001010000011" & 
    "0010001011010010" & 
    "1110000010101100" & 
    "0000101101111011" & 
    "1101111100000101" & 
    "1111111110101100" & 
    "0000010001000000" & 
    "1100110100010101" & 
    "1111111110110110" & 
    "1110011110101010" & 
    "0001101011011111" & 
    "0010101111110111" & 
    "1111100101111101" & 
    "0010000111110001" & 
    "1111100011001001" & 
    "1110100111101011" & 
    "1111110001101101" & 
    "1101011100100111" & 
    "0001101101010001" & 
    "1110101110111001" & 
    "0010000000100000" & 
    "0000011010110111" & 
    "0000101010000010" & 
    "0001111011111111" & 
    "1110000010111010" & 
    "1111110111001110" & 
    "0000111111000000" & 
    "1110101101011101" & 
    "1111000100101000" & 
    "1101100100101001" & 
    "1111101000001111" & 
    "1110101011011011" & 
    "1111111110101000" & 
    "0000101010110001" & 
    "0001101110101001" & 
    "0000001100101010" & 
    "0001011110100001" & 
    "1110011001100010" & 
    "0000100101011110" & 
    "1110011010010001" & 
    "0000000100101011" & 
    "0000010100100100" & 
    "1110011111111101" & 
    "1111110100010110" & 
    "1111100101001011" & 
    "0001001010111011" & 
    "0000111101110001" & 
    "0000101000110111" & 
    "0010011010011011" & 
    "1111000101001001" & 
    "0001100110101100" & 
    "1111101101101111" & 
    "1110001010010101" & 
    "0000010111100011" & 
    "1101111001000011" & 
    "1111001111110101" & 
    "0000010001000101" & 
    "0000000011001111" & 
    "0001000111000111" & 
    "0000001111110110" & 
    "0001000010100001" & 
    "0001100000011101" & 
    "0000010111000010" & 
    "0000101100010011" & 
    "1111010001110100" & 
    "0000010001011101" & 
    "1111011110001011" & 
    "1111111011011100" & 
    "1111100101010010" & 
    "1110000001110011" & 
    "1110100111110011" & 
    "0001110000010110" & 
    "0000111011110011" & 
    "0001111010111001" & 
    "0000111101110100" & 
    "0001000001110101" & 
    "0000101010011010" & 
    "1110111000001101" & 
    "0000101000011000" & 
    "1110010011001111" & 
    "0010001010101010" & 
    "1110100000010100" & 
    "1101001001100100" & 
    "0000001010110010" & 
    "1110110100111010" & 
    "0000110110000001" & 
    "0001000110111111" & 
    "1111101100111001" & 
    "0001110110011011" & 
    "1111011001001001" & 
    "0000011011000100" & 
    "0001001010000101" & 
    "1111011011000000" & 
    "1110111010000110" & 
    "1100011011111011" & 
    "0001010001100001" & 
    "1111000000100110" & 
    "0000001000100101" & 
    "0010000010010001" & 
    "0010010010110110" & 
    "0000110001101001" & 
    "1111110111010101" & 
    "1111000000000100" & 
    "0000011011111101" & 
    "1110010001001101" & 
    "1110110001010101" & 
    "1110011100101111" & 
    "1111010100011111" & 
    "1111111101110101" & 
    "1110111000110100" & 
    "0010100110111110" & 
    "0000110110111101" & 
    "1111110001111001" & 
    "0010001101010111" & 
    "1110101101000001" & 
    "0000101100110111" & 
    "1111000010001100" & 
    "1111001101100011" & 
    "0000110100100000" & 
    "1110100011010110" & 
    "1111100000011001" & 
    "1111110011010100" & 
    "1111110011000001" & 
    "0001100011111101" & 
    "1111101010001010" & 
    "0001110101000001" & 
    "0000000100110000" & 
    "1111111010001011" & 
    "1111101010001101" & 
    "1111001010111110" & 
    "1110110110110110" & 
    "1111110110010010" & 
    "1111111110010111" & 
    "0000111001010010" & 
    "1111011110110101" & 
    "0011010001111111" & 
    "0010001110101000" & 
    "1111011111001111" & 
    "0001111101010100" & 
    "1110101001001100" & 
    "0000011000001010" & 
    "0000110010111001" & 
    "1100100110000010" & 
    "0001001110000100" & 
    "0000001110010010" & 
    "0000011010110101" & 
    "0010100101110101" & 
    "0000001110010000" & 
    "0000110000110101" & 
    "1101110111111011" & 
    "0000100000101111" & 
    "0001000101011110" & 
    "1111000101010010" & 
    "0000100110101100" & 
    "1101100111110011" & 
    "1111100001011111" & 
    "1110000010000111" & 
    "1110001111100101" & 
    "0000011111011000" & 
    "0000011100001001" & 
    "0001010000110111" & 
    "0000000111110100" & 
    "1111111010010001" & 
    "0000100111101000" & 
    "1110010101100100" & 
    "0000100010010010" & 
    "1111011111100010" & 
    "1110100110001110" & 
    "0001000100110011" & 
    "1110111100100001" & 
    "0000111011000011" & 
    "0001100001110010" & 
    "0001001111001110" & 
    "0010011110011101" & 
    "0001011110101100" & 
    "0000110111100001" & 
    "0000010100101111" & 
    "0000011101110111" & 
    "1111101011100110" & 
    "1110001100100011" & 
    "0000010011001001" & 
    "1111110100100100" & 
    "0000011010001001" & 
    "0010010101111101" & 
    "0000001101100010" & 
    "0000100000000000" & 
    "0001110110000010" & 
    "1110100010011001" & 
    "0001100011011011" & 
    "1111110011111110" & 
    "1111111000100111" & 
    "0000010000100101" & 
    "0000001111001110" & 
    "0001000111010111" & 
    "1111000010000100" & 
    "0001000000110111" & 
    "0001010001010011" & 
    "1110110000001011" & 
    "0001100101010110" & 
    "0001010010101100" & 
    "0000110011010010" & 
    "0000111101000101" & 
    "1101110000100100" & 
    "0000010000010111" & 
    "1110110011001001" & 
    "1110000001001001" & 
    "0000000001001111" & 
    "1110110100100110" & 
    "0000010111101001" & 
    "1111111000011110" & 
    "1111011000011010" & 
    "1111001001100101" & 
    "1110101111100011" & 
    "0000010100011001" & 
    "1101110101001010" & 
    "1101111100100011" & 
    "1111101010101110" & 
    "1100100110101101" & 
    "0000010011010010" & 
    "1111100011010110" & 
    "0000010111101010" & 
    "0000111100000010" & 
    "1111101100000111" & 
    "0000100001000111" & 
    "0000000001100000" & 
    "0001110011100100" & 
    "0010000111000011" & 
    "1110010101011100" & 
    "1110100100000101" & 
    "1110010111011000" & 
    "1111110000010111" & 
    "1111011100011101" & 
    "1101110110101101" & 
    "0011010101010101" & 
    "1101100011111000" & 
    "0000110001001000" & 
    "1111111101001100" & 
    "1111010010001011" & 
    "0001101000001000" & 
    "1111001001000100" & 
    "1110111101100000" & 
    "0000001010000000" & 
    "1110110100100100" & 
    "0000110101101010" & 
    "1110010101101111" & 
    "0001011010111010" & 
    "0001100000010111" & 
    "0010100100111000" & 
    "0011000100000100" & 
    "0001001110010110" & 
    "0000111001011101" & 
    "1111000101010110" & 
    "1110011001001110" & 
    "1111011011101110" & 
    "1101101000101001" & 
    "1111111011110011" & 
    "1111000111010110" & 
    "1110000110111100" & 
    "0000111001100101" & 
    "1111110000100101" & 
    "0001101011111110" & 
    "0000010100110011" & 
    "0000001111001100" & 
    "0001011000110001" & 
    "0000010100111111" & 
    "1111011101010110" & 
    "1111001111101011" & 
    "1101000001110001" & 
    "1110110011100100" & 
    "1111000100110110" & 
    "0000000111110101" & 
    "0001010110010100" & 
    "1111001011001011" & 
    "0011111010001001" & 
    "0000001100001000" & 
    "0001111001000101" & 
    "0000001001010001" & 
    "1110100110100101" & 
    "0000111000011001" & 
    "1110110000010011" & 
    "1110010000100101" & 
    "1110001000111001" & 
    "1101111001111110" & 
    "1111111001001011" & 
    "1111111110101100" & 
    "0000110111011101" & 
    "0000111010001110" & 
    "1110100011110010" & 
    "0010000101101011" & 
    "1111011100010111" & 
    "1111100101010000" & 
    "0000011001101000" & 
    "1101010100110011" & 
    "0000100110110001" & 
    "1111000111010001" & 
    "0000101110001001" & 
    "0000000111011001" & 
    "0000011001001110" & 
    "0001011111000011" & 
    "1111001010111100" & 
    "1111101001000100" & 
    "0001011010001110" & 
    "1101111010110101" & 
    "0000000001001010" & 
    "1100111111011000" & 
    "1111000101010000" & 
    "1100011100001000" & 
    "1101111010101011" & 
    "1111111000011111" & 
    "1110111001111101" & 
    "0001000100001000" & 
    "0000111100111100" & 
    "0001110111010100" & 
    "0000101111001100" & 
    "1110110000001111" & 
    "1110000110100011" & 
    "1110111001101110" & 
    "1100110111000110" & 
    "0000001110001010" & 
    "1111100111100101" & 
    "0000110001101011" & 
    "0000001001001111" & 
    "1110011011111101" & 
    "0011011101011100" & 
    "0010000111100001" & 
    "0000111101110010" & 
    "1111011000011100" & 
    "1111111101101000" & 
    "1111100110010011" & 
    "1101101110101010" & 
    "0000010001000000" & 
    "1110010010010101" & 
    "1101000011000000" & 
    "0001101110101101" & 
    "0000010100100010" & 
    "0001010111110111" & 
    "0001110001100011" & 
    "0001000000001001" & 
    "0010010001111001" & 
    "1110011011110110" & 
    "0000011110110100" & 
    "1111100011010111" & 
    "1101101100011000" & 
    "1110111111110110" & 
    "1111011010011000" & 
    "0000000001001010" & 
    "0000111001000011" & 
    "1111010001100100" & 
    "0000011100110001" & 
    "0000001111010010" & 
    "0000110010000110" & 
    "0001100100100010" & 
    "1111100100010010" & 
    "0001001111101001" & 
    "1101011100110011" & 
    "1110011100010110" & 
    "1110011001110001" & 
    "1111100000000110" & 
    "0100000110010010" & 
    "0000101001011100" & 
    "0000100000010011" & 
    "0010000111010100" & 
    "1110110010101010" & 
    "1111111000100111" & 
    "1111101110001001" & 
    "1110111001001101" & 
    "1111101100100000" & 
    "1111100110110000" & 
    "0000100101111001" & 
    "1111101100011110" & 
    "1110110001000010" & 
    "0001100000011010" & 
    "0010001101001011" & 
    "0010100010101001" & 
    "1110100001101100" & 
    "0000101001000100" & 
    "1111110111110011" & 
    "1111001001011111" & 
    "0000100110100110" & 
    "1110100110101011" & 
    "1111000000111111" & 
    "1111000100101000" & 
    "1110011010100000" & 
    "0010001010011010" & 
    "1110000100010010" & 
    "0001000100100000" & 
    "0001100011000101" & 
    "1111010001000110" & 
    "0001110010010100" & 
    "1110111011101011" & 
    "1110101110111100" & 
    "1111100010100110" & 
    "1101111011100100" & 
    "1111110001111111" & 
    "1110000011011101" & 
    "0000011011101111" & 
    "1110111111111011" & 
    "1111101010110100" & 
    "0001011101001110" & 
    "1111001001111100" & 
    "0001011111110110" & 
    "1111101000110011" & 
    "1111010011100101" & 
    "0001001010101011" & 
    "1110000010101100" & 
    "1111101010000011" & 
    "0000010011111010" & 
    "1110111011000011" & 
    "0001110110011001" & 
    "1110101010000101" & 
    "0010011000110101" & 
    "0000010010011100" & 
    "1110000101110101" & 
    "0010101100011001" & 
    "1110111100001110" & 
    "0000000111101110" & 
    "1111000001000001" & 
    "1101001011011010" & 
    "1101000111100011" & 
    "1111011001000100" & 
    "0000000101011101" & 
    "0000101001011100" & 
    "0000011110010001" & 
    "0000100101001010" & 
    "1111010101101000" & 
    "0001111111100000" & 
    "0000111110000100" & 
    "1101011110111110" & 
    "1101111111001110" & 
    "1101101000001011" & 
    "1111100101111110" & 
    "0000100111010011" & 
    "1111000110001111" & 
    "0000001011111101" & 
    "0000001110011110" & 
    "0000000110101111" & 
    "0000010100010001" & 
    "1111010001000010" & 
    "0000000101000110" & 
    "1110101110111001" & 
    "1110110001011001" & 
    "1111000101111111" & 
    "1101101111001000" & 
    "1111110010000000" & 
    "1110010000110000" & 
    "0001100110101111" & 
    "0001011101001000" & 
    "0000001000000110" & 
    "0000100010000111" & 
    "1110011100010000" & 
    "1110111000010101" & 
    "0010111110100010" & 
    "1111101111001101" & 
    "0000011100101011" & 
    "1101001110011000" & 
    "1110001110111010" & 
    "0000001110000010" & 
    "0000100100011001" & 
    "1111100111011010" & 
    "1111011110000111" & 
    "0001001100011000" & 
    "1111010010010010" & 
    "0000110000101110" & 
    "0000111001001111" & 
    "0000111010100111" & 
    "1111010001111110" & 
    "1111110010011101" & 
    "1101000011100111" & 
    "1111100100001111" & 
    "1101100110001011" & 
    "0000110000111011" & 
    "0010001001011001" & 
    "1111011110010100" & 
    "0010011011111011" & 
    "1111100100000010" & 
    "0000111100100111" & 
    "0001100100010111" & 
    "1110111000101011" & 
    "1111001001110111" & 
    "1101010101111000" & 
    "1111001101011010" & 
    "1111011110101110" & 
    "1110001000110100" & 
    "0001011111010110" & 
    "0001001011111100" & 
    "0001000001101100" & 
    "0001000100101011" & 
    "1101101101111111" & 
    "0000100010001101" & 
    "1101100111000100" & 
    "1111010010010001" & 
    "1111111001111010" & 
    "1111101110001110" & 
    "0001111111010101" & 
    "1110101001100000" & 
    "0000000011010011" & 
    "0001101010011001" & 
    "0000100011101011" & 
    "0010110000111110" & 
    "0000110110000111" & 
    "1111010111010101" & 
    "0000111010011000" & 
    "1110101011000111" & 
    "1111011011100100" & 
    "1101100000010110" & 
    "0000101010010010" & 
    "1110110111001010" & 
    "1101110001000101" & 
    "0001100001100001" & 
    "0001111011100100" & 
    "0001010011011010" & 
    "0001100101100000" & 
    "1110111110110101" & 
    "0010111110111011" & 
    "1111001000001111" & 
    "0000001100111010" & 
    "1110011011010110" & 
    "1111000011011001" & 
    "0000100101001000" & 
    "1101100110111111" & 
    "0000011010010110" & 
    "0000011001001111" & 
    "0000001011010011" & 
    "0001101111111110" & 
    "1111111000001010" & 
    "1111110011111110" & 
    "0000000011000111" & 
    "1111100010000010" & 
    "0001111011111000" & 
    "1101000010011101" & 
    "0001110000011011" & 
    "0001001100101010" & 
    "1111001011000001" & 
    "0001000000100000" & 
    "1111001110001010" & 
    "0010000111000100" & 
    "0000100101010100" & 
    "1111011101010100" & 
    "0010001100010101" & 
    "1111011100001000" & 
    "0000100100011000" & 
    "1111111000100101" & 
    "1101110011000100" & 
    "1111101011010110" & 
    "1111100011111100" & 
    "1111101100110110" & 
    "0010000010000001" & 
    "0000110110111010" & 
    "0010010010011011" & 
    "0000000100100001" & 
    "0001001101011110" & 
    "0011111001100000" & 
    "1110101001110010" & 
    "1110101000100110" & 
    "0000000111010011" & 
    "1111111111010011" & 
    "1111000001100001" & 
    "0001100111101111" & 
    "0001110111000010" & 
    "0000001101101101" & 
    "0000011111111111" & 
    "0000001101100111" & 
    "1110001001101101" & 
    "0000111000101101" & 
    "1101111100110101" & 
    "0000010100011100" & 
    "1111000011111100" & 
    "1111111101111100" & 
    "0001101100111010" & 
    "1110111011011110" & 
    "0000000101101101" & 
    "0001111111110100" & 
    "1110111010111100" & 
    "0010101011000111" & 
    "1111011001011111" & 
    "0000011100011101" & 
    "1111101100110011" & 
    "1111010101110100" & 
    "1111011010011011" & 
    "1101001000101010" & 
    "1111111011101010" & 
    "1111001111111000" & 
    "1111010111011000" & 
    "0000111101010000" & 
    "0000001100001000" & 
    "1110101101101001" & 
    "0001101111100101" & 
    "0001110001100000" & 
    "0010010110010011" & 
    "1111111010100010" & 
    "1111011011101001" & 
    "1111100011110111" & 
    "1110011100010111" & 
    "0000010010011001" & 
    "1101111011110101" & 
    "0000000001010000" & 
    "0000101010111001" & 
    "1111100101100011" & 
    "0010110101100100" & 
    "0010100110110001" & 
    "1111100001011000" & 
    "0000100000000001" & 
    "1101010100101010" & 
    "0001011111100101" & 
    "1111100110111110" & 
    "1101101101111000" & 
    "0001100111011000" & 
    "1101111010110100" & 
    "0001100010010011" & 
    "0001000001001101" & 
    "0001011011001100" & 
    "0011100100101100" & 
    "0010101011000011" & 
    "0001011100101000" & 
    "1101000110001011" & 
    "1111010011101000" & 
    "1110100010000000" & 
    "1101011011110010" & 
    "1111000100000011" & 
    "1110110101111111" & 
    "0010011110101000" & 
    "0000001000010000" & 
    "1111110010010111" & 
    "0011001010101010" & 
    "0001010001111011" & 
    "0001010101001001" & 
    "0001011001011101" & 
    "1111101000101101" & 
    "1111110011110011" & 
    "1110101000001011" & 
    "1111000101001000" & 
    "1110110001011001" & 
    "1111101000110111" & 
    "0001011000000110" & 
    "1111101110111010" & 
    "0001100100011100" & 
    "0010010000111111" & 
    "0000010100000010" & 
    "0001100000001111" & 
    "1111010010001001" & 
    "1111101110010001" & 
    "1110100110101101" & 
    "1110111111000101" & 
    "0001100110011001" & 
    "1110001110110011" & 
    "0010010011001011" & 
    "0000101010110011" & 
    "1111110100101101" & 
    "0001000110100011" & 
    "1111010001100110" & 
    "1111111001000101" & 
    "0000101110011101" & 
    "0000010111001100" & 
    "0000101101111111" & 
    "1111000011011001" & 
    "0000101110001010" & 
    "1101001011000001" & 
    "1110110101100000" & 
    "0001101010011000" & 
    "0000101000110010" & 
    "1111111110010000" & 
    "0000010001011001" & 
    "0000101101011111" & 
    "0001001100010100" & 
    "1111100011101000" & 
    "1110101101100000" & 
    "1101101111101101" & 
    "1110111101011100" & 
    "0001011000100110" & 
    "0000011001011011" & 
    "1110110101101111" & 
    "1111100000100001" & 
    "1110100101111111" & 
    "0001111101010101" & 
    "1111011100111011" & 
    "0010001010001011" & 
    "1110111010101011" & 
    "1101000001011110" & 
    "0000011001010111" & 
    "1111011001000101" & 
    "1110100100111001" & 
    "1110011001111111" & 
    "1110110110101011" & 
    "1111101011000011" & 
    "1111111011111111" & 
    "0010000110110010" & 
    "0001011111101101" & 
    "1110000000101100" & 
    "0000110001011011" & 
    "1110101100111010" & 
    "0001011111000011" & 
    "0000010010110101" & 
    "1110001001000101" & 
    "0001100000000001" & 
    "1101101110000111" & 
    "0000000001100000" & 
    "0010010000011110" & 
    "0001100100011101" & 
    "0010101110110000" & 
    "0000100011101110" & 
    "0000010000100100" & 
    "0001000111011110" & 
    "1101111011111110" & 
    "0000110001000000" & 
    "1110011110110001" & 
    "0000100001001100" & 
    "1111001111101110" & 
    "1111101000111100" & 
    "0010000110100011" & 
    "1111000001011000" & 
    "0001011011110001" & 
    "0010110111111111" & 
    "0000000010000101" & 
    "0001000000000010" & 
    "1111011101011101" & 
    "1111011001011000" & 
    "1111110100101000" & 
    "1110000100000111" & 
    "0000001011000011" & 
    "1111001110011110" & 
    "0001101110111111" & 
    "0001010010111111" & 
    "0001101101110011" & 
    "1111111110001100" & 
    "1111100111100011" & 
    "0001000101001011" & 
    "1111100010010110" & 
    "1101011111010100" & 
    "0000110011101110" & 
    "1110110011111100" & 
    "1111101010110011" & 
    "0000000100010010" & 
    "1110001000100001" & 
    "0000110011111011" & 
    "1111110100000011" & 
    "0000100101110000" & 
    "0001100111000000" & 
    "0010010010010000" & 
    "0000110100111011" & 
    "1111101001101011" & 
    "1110101000110010" & 
    "0000101110000000" & 
    "1101001110101101" & 
    "0000011001100101" & 
    "1110001001011001" & 
    "0000111000100100" & 
    "0000110110110011" & 
    "0000000001011111" & 
    "0100111100101111" & 
    "1111011011111111" & 
    "0000110011000100" & 
    "0011000011100001" & 
    "1101100111100101" & 
    "0000101111100111" & 
    "1101000111110101" & 
    "0000011010001111" & 
    "1111111111111100" & 
    "1111101001111110" & 
    "0001000001111100" & 
    "0000001010100100" & 
    "0010110000000000" & 
    "1111000000001010" & 
    "1110010010010110" & 
    "0001101110010111" & 
    "1110010110010101" & 
    "1111011000000001" & 
    "1101111000011110" & 
    "1101010010110100" & 
    "1111110010010111" & 
    "1110000010100001" & 
    "1111100000010110" & 
    "0000011011000101" & 
    "1111000111111110" & 
    "0011010101111000" & 
    "1111000101000011" & 
    "0010101010011011" & 
    "1111111111110101" & 
    "1101010100000100" & 
    "1111100100101000" & 
    "1111001000100010" & 
    "0000011011110110" & 
    "1111110101001111" & 
    "1111010010101000" & 
    "0001111100010010" & 
    "1110011101100000" & 
    "0000101100100010" & 
    "1111011100101001" & 
    "1111011110001001" & 
    "0010010000100010" & 
    "1111101110001001" & 
    "0001111101011010" & 
    "1111100010111100" & 
    "1100000010101110" & 
    "0001111000010110" & 
    "0000000011000010" & 
    "1111110010100000" & 
    "0001000100010100" & 
    "0000110110001100" & 
    "0010011000101000" & 
    "0000110000111000" & 
    "0000101110110111" & 
    "0000010101010100" & 
    "1110110110100111" & 
    "1111011001101100" & 
    "1111100111110011" & 
    "1111011000101011" & 
    "0000010110111011" & 
    "1110001001100001" & 
    "0000001110111110" & 
    "1111110101000100" & 
    "0001000001100110" & 
    "0010011110001111" & 
    "0000100001101011" & 
    "0001110110011000" & 
    "1101100011110000" & 
    "1110101101000011" & 
    "1111100101001101" & 
    "1101110110011110" & 
    "0001011110110010" & 
    "0000000110110100" & 
    "1111110010101000" & 
    "0001101110000101" & 
    "0001011101100111" & 
    "0010010100100011" & 
    "0001101100001101" & 
    "0001111010000100" & 
    "0000100101100000" & 
    "1111101001000110" & 
    "0000011000101011" & 
    "1101110010001011" & 
    "1111101111001110" & 
    "1111101101010011" & 
    "1110101000111001" & 
    "0011000101001000" & 
    "0000001001000010" & 
    "0100000000100001" & 
    "0000111110110100" & 
    "0000011110111111" & 
    "0010111001000100" & 
    "0001101110111010" & 
    "1111111110011010" & 
    "1110100101101100" & 
    "1111000000001001" & 
    "1110110111110000" & 
    "1110011111011101" & 
    "0000101001001100" & 
    "0010010101011010" & 
    "0001100000010010" & 
    "0001111110001111" & 
    "0000111111011100" & 
    "0000100001100001" & 
    "0001000010000111" & 
    "0000101011100011" & 
    "0000010110010000" & 
    "1101111001100000" & 
    "1110111000010001" & 
    "0000011000110110" & 
    "0000010101110100" & 
    "0011011011110101" & 
    "1111111110010101" & 
    "0001011100001101" & 
    "0000101001010001" & 
    "0001100010000011" & 
    "0001001110111101" & 
    "1110100001111100" & 
    "0001110110110001" & 
    "0000001100000111" & 
    "1110111010100101" & 
    "1111001011110111" & 
    "1111001100110000" & 
    "0000111001000101" & 
    "1111110000001011" & 
    "1111110101110111" & 
    "0001100110000101" & 
    "0000100110000110" & 
    "1111110101101000" & 
    "0001011101100000" & 
    "0000100011001101" & 
    "1111111000110010" & 
    "1110001100001011" & 
    "1111111000101101" & 
    "0000110111111111" & 
    "1111100001101001" & 
    "0001101101001100" & 
    "1111011011111111" & 
    "0001000010111101" & 
    "0001111001000001" & 
    "0001100110100101" & 
    "0001111000001010" & 
    "1101110011000011" & 
    "0000000110101101" & 
    "1111010010011000" & 
    "1101111101000111" & 
    "1111111110001100" & 
    "1101111000101011" & 
    "0000000011010001" & 
    "0000000011111000" & 
    "1111101100111101" & 
    "0010000111100000" & 
    "0000001111011110" & 
    "0000101000010001" & 
    "0000001110000010" & 
    "1110110011001000" & 
    "0000101001100011" & 
    "1111011110110000" & 
    "1111111111111101" & 
    "1111011000101001" & 
    "1111100110100000" & 
    "0001000100000100" & 
    "1110001000111010" & 
    "1110111011100011" & 
    "1111100100000110" & 
    "1111101011101101" & 
    "0000101100001000" & 
    "1110010010001001" & 
    "1111101101100101" & 
    "1110101110000110" & 
    "1101100100011000" & 
    "0000110011001111" & 
    "1111100011000011" & 
    "0010110011101111" & 
    "0001001001011011" & 
    "0000001000000010" & 
    "0001011011010000" & 
    "1111110111110100" & 
    "0000110010110110" & 
    "1110100111011011" & 
    "1110100000100000" & 
    "0000111100001100" & 
    "1101101000001101" & 
    "1111110111111010" & 
    "0000101010011100" & 
    "0000000101001011" & 
    "0010000101100000" & 
    "1101101010010000" & 
    "0000101101101001" & 
    "0010001011011110" & 
    "0000010100001001" & 
    "0001010100000110" & 
    "1111011100001100" & 
    "0000110011010100" & 
    "1111100010000111" & 
    "1101011100001011" & 
    "0000000000101100" & 
    "1110100011101011" & 
    "0001010001001100" & 
    "0001010000011101" & 
    "0000100111010110" & 
    "0010001001011110" & 
    "1111101101001000" & 
    "0000111001111111" & 
    "0000100101101011" & 
    "1101010111100000" & 
    "0000010111101011" & 
    "1111001000000110" & 
    "1111010001001110" & 
    "0001001111100111" & 
    "1111100100000111" & 
    "0000111000111000" & 
    "1111110001000010" & 
    "0001000000001010" & 
    "0001100001001101" & 
    "0000101011001011" & 
    "0001000001000110" & 
    "1111011101100101" & 
    "0001011011010101" & 
    "0000010011111001" & 
    "1111000001100011" & 
    "1111011000000101" & 
    "1110001110110010" & 
    "0000100111010100" & 
    "0000101111101000" & 
    "1110011100010011" & 
    "0000011111000101" & 
    "0001000101111111" & 
    "0000000101100011" & 
    "0010011100110100" & 
    "1100100010110001" & 
    "0000101000111100" & 
    "1110001100110001" & 
    "1110100111111000" & 
    "0000000100110111" & 
    "1110001101011011" & 
    "0010001010110011" & 
    "1111111111001010" & 
    "1111101000110110" & 
    "1110110110100101" & 
    "1111101000101110" & 
    "0010011101000111" & 
    "1111001011110101" & 
    "1111101110011101" & 
    "0000000100010010" & 
    "1100110011100011" & 
    "0001100111011101" & 
    "1101110111110001" & 
    "0000011010001110" & 
    "0000011110110011" & 
    "0000001101111000" & 
    "0000000011100011" & 
    "0001100101110101" & 
    "0001011001000000" & 
    "0010011000011100" & 
    "0000001011101001" & 
    "0000001100111101" & 
    "1101010000101000" & 
    "1101101000111111" & 
    "1111101100000100" & 
    "1111001110010000" & 
    "0010010110101101" & 
    "1110111110000001" & 
    "0010000100101001" & 
    "0001010110010110" & 
    "1111001001010111" & 
    "0010000101010101" & 
    "1111010001001111" & 
    "1111011011111100" & 
    "0001010000011011" & 
    "1110110011101110" & 
    "0000000101001011" & 
    "1111000010101111" & 
    "0000011101010111" & 
    "0001000001001100" & 
    "0000100001010110" & 
    "0001011001011000" & 
    "1111010001010011" & 
    "0001001101001010" & 
    "0010010000011100" & 
    "1110011101010110" & 
    "1111001011011010" & 
    "1101111101011101" & 
    "1110111001010011" & 
    "1111010110000010" & 
    "1111011110101010" & 
    "0001001011011101" & 
    "1111010100110110" & 
    "0000110101010111" & 
    "1111111101001000" & 
    "1111000011111000" & 
    "1111111001010110" & 
    "1110011111001101" & 
    "1110100101100010" & 
    "1110101011000001" & 
    "1101111001011011" & 
    "1110111111011001" & 
    "1110101111101111" & 
    "0000101101100101" & 
    "1111111000011011" & 
    "0001001011100110" & 
    "0000011010011111" & 
    "1111101011001111" & 
    "1111010111000011" & 
    "0000000001101111" & 
    "1101011100010000" & 
    "1111100111011100" & 
    "1101011101010101" & 
    "1110001100011100" & 
    "1101100110110101" & 
    "1111100100011001" & 
    "0011010011110010" & 
    "0010001001001011" & 
    "0000110010010001" & 
    "0001001110110101" & 
    "1111011101000100" & 
    "0001011000101001" & 
    "1110000101011011" & 
    "1101110000001001" & 
    "1111010101111100" & 
    "1100111110010100" & 
    "1110010010011110" & 
    "0001001000111011" & 
    "0000001000110111" & 
    "0001001111111011" & 
    "0001010000101000" & 
    "0000010100001011" & 
    "0000011110110000" & 
    "0001010110001100" & 
    "0000011101000111" & 
    "1110111011000101" & 
    "1111101010011100" & 
    "1110111011000000" & 
    "1110100001111000" & 
    "1110111000000001" & 
    "1111101110101010" & 
    "0010111111101110" & 
    "1111100010001001" & 
    "0000110001011100" & 
    "0001101011111001" & 
    "0000111111100000" & 
    "0010010001101111" & 
    "1111010001100001" & 
    "1111000010011000" & 
    "0000000000100101" & 
    "1110000111101010" & 
    "0001100100010110" & 
    "1101010110110110" & 
    "0000100000110101" & 
    "0010001000100111" & 
    "1111100100101000" & 
    "0001011000000001" & 
    "1111001000100011" & 
    "0000100100001111" & 
    "0000001010111110" & 
    "1110111001101110" & 
    "1111010011101100" & 
    "1110010010000001" & 
    "1110110001101000" & 
    "1111010011011001" & 
    "1110001010100110" & 
    "0001000001101101" & 
    "0011011111010110" & 
    "0100101011110110" & 
    "0010011011001011" & 
    "0000101101010001" & 
    "0000000001111110" & 
    "1110011010110100" & 
    "1111000011010110" & 
    "1111111010100010" & 
    "1110101011101001" & 
    "0000010011001011" & 
    "1110011011001100" & 
    "1111011100100011" & 
    "0000110110011010" & 
    "0001001101001110" & 
    "0010011011010110" & 
    "0000001111111001" & 
    "0001100000001010" & 
    "0000111101001100" & 
    "1101001001100001" & 
    "0000001101011011" & 
    "1101110001011110" & 
    "1101010110000110" & 
    "1110010101111101" & 
    "1110101011110001" & 
    "0010001000100111" & 
    "1111101100001101" & 
    "0001100010100011" & 
    "0000011000010011" & 
    "1101110000110100" & 
    "0001011001110010" & 
    "1110000011010111" & 
    "0000110110000010" & 
    "0001000111010100" & 
    "1101110100111100" & 
    "0001011000100100" & 
    "1111101110000000" & 
    "1110111101001111" & 
    "0000110011111100" & 
    "0000010101000001" & 
    "0010100001011110" & 
    "0000101111101000" & 
    "0001100001001111" & 
    "0001000011001110" & 
    "1110011100111110" & 
    "0000100100100000" & 
    "1011111100100011" & 
    "1110001101100000" & 
    "0000110111111010" & 
    "1110010101111100" & 
    "0001101000101111" & 
    "0001011011011001" & 
    "0000011000111000" & 
    "0000010100011000" & 
    "1111011011010110" & 
    "0001110000000000" & 
    "1110110011001000" & 
    "1110101100011010" & 
    "1101110011100111" & 
    "1101110101000010" & 
    "1111111110000100" & 
    "1110001110101110" & 
    "0000000111000010" & 
    "1111101111111110" & 
    "0000100111011101" & 
    "1111110100110101" & 
    "0000001101100100" & 
    "0001100000111001" & 
    "1111100001011110" & 
    "1110101101010100" & 
    "0000011110111001" & 
    "1101100101011001" & 
    "1111010111011001" & 
    "0000000101010111" & 
    "1110000100010000" & 
    "0010001001001111" & 
    "0001000000111011" & 
    "0001100110010101" & 
    "0001010010101111" & 
    "1110110000010110" & 
    "0001110011011101" & 
    "1101110010011011" & 
    "0001010000110011" & 
    "1111111001111110" & 
    "1110011101101011" & 
    "1111110011000010" & 
    "1100100101101100" & 
    "1111001011010010" & 
    "0001001101011101" & 
    "0010011110101101" & 
    "0010101111011000" & 
    "0000011000001000" & 
    "0000010011011001" & 
    "0000011111101000" & 
    "1111101110100100" & 
    "1111111011111110" & 
    "0000000101110011" & 
    "1110001010001011" & 
    "1111010010111010" & 
    "1111000011100110" & 
    "1111010110101110" & 
    "0000011111000100" & 
    "0001010110110000" & 
    "0001010110111100" & 
    "0000101101101111" & 
    "0010010110100101" & 
    "1111110011100101" & 
    "1111001100111111" & 
    "1111010101010011" & 
    "1110100011010110" & 
    "1110111011110010" & 
    "1101101110101011" & 
    "1111111100011110" & 
    "0000111011000011" & 
    "0001110110111011" & 
    "0010110011000010" & 
    "1111100111111111" & 
    "0000001101110100" & 
    "0001111001111101" & 
    "0001011111111011" & 
    "0000010110111100" & 
    "1101101110000101" & 
    "1101111101110111" & 
    "0000101001011000" & 
    "1111010010110001" & 
    "0010011110010111" & 
    "1111000000101110" & 
    "0001100001001010" & 
    "0000100111111010" & 
    "0001001100011110" & 
    "0000110000100000" & 
    "1110111010101001" & 
    "1111010100101110" & 
    "0000010111111001" & 
    "1110101000001001" & 
    "1111001011111101" & 
    "1110001000011111" & 
    "1111010100111000" & 
    "0001010110011100" & 
    "0000011001100011" & 
    "0000010111010101" & 
    "1110001010010001" & 
    "0000110011011111" & 
    "0001000100011011" & 
    "1110111011110010" & 
    "1110101001011011" & 
    "1100101001011010" & 
    "0000001111110001" & 
    "1111100001101011" & 
    "1110100111100001" & 
    "0010101000000001" & 
    "1111000111111010" & 
    "0001011010011100" & 
    "0001101100100000" & 
    "0000101111010110" & 
    "0000011101000110" & 
    "1111010111000110" & 
    "0010011010111001" & 
    "1101110111011100" & 
    "1110101000100000" & 
    "1111111101100001" & 
    "1101111100000011" & 
    "1111100010100011" & 
    "0001010101111100" & 
    "0010011000100000" & 
    "0001001101001100" & 
    "0000100110111011" & 
    "0000010010010011" & 
    "0010010110010011" & 
    "1111010011110101" & 
    "0000000011011001" & 
    "1110110100011010" & 
    "1111010111111011" & 
    "0000110001110110" & 
    "1110110100010111" & 
    "0000001100000000" & 
    "0000001010101010" & 
    "0010110101101011" & 
    "0000000101001100" & 
    "1111101011010111" & 
    "0010010100000110" & 
    "1101000101010110" & 
    "0000010011000001" & 
    "0000001000011101" & 
    "1110011010011001" & 
    "1111011010111011" & 
    "1110110000100001" & 
    "0000011101110001" & 
    "0001110001111011" & 
    "0000101110110001" & 
    "0001101001100101" & 
    "0001101011111111" & 
    "0000110010110100" & 
    "1111100011110010" & 
    "1110010100111011" & 
    "0001000011001011" & 
    "1110011001001110" & 
    "0000010001001010" & 
    "1111101111011010" & 
    "0001011111011001" & 
    "1111101001001011" & 
    "1111100000010000" & 
    "0001001100011000" & 
    "0001010111011111" & 
    "0001011000000101" & 
    "0001100001110101" & 
    "1110111000111000" & 
    "1111101111011000" & 
    "0000001000010111" & 
    "1101100000100111" & 
    "0000101001000101" & 
    "1101001100110100" & 
    "0000010010110000" & 
    "1111111001110011" & 
    "1111011010100001" & 
    "0010010010000101" & 
    "1110111100010011" & 
    "1111110110110010" & 
    "1110110110110010" & 
    "1100100010010110" & 
    "0000000010100010" & 
    "1111010111001001" & 
    "1111001100101000" & 
    "1111011100000001" & 
    "1101111101001111" & 
    "0010111001000111" & 
    "1111101010111011" & 
    "0010100100100101" & 
    "0001101000111100" & 
    "1111101010000011" & 
    "0010011001000010" & 
    "1111111111000111" & 
    "1111100011110110" & 
    "0000101011001110" & 
    "1111111110101111" & 
    "0000001000000010" & 
    "1110100000100111" & 
    "0000110001101100" & 
    "0001001100100101" & 
    "0000110111111111" & 
    "0001101111101001" & 
    "0000110010000101" & 
    "0001111001001100" & 
    "0000100011001010" & 
    "1110111010110010" & 
    "1110111011111101" & 
    "1101000001101011" & 
    "1101111010101111" & 
    "1110011011010110" & 
    "1110110110010011" & 
    "1111101100011011" & 
    "0010001010101000" & 
    "0010000001000101" & 
    "1111001101011100" & 
    "1110110000111111" & 
    "0001001100111011" & 
    "1101010010100111" & 
    "1111001101100011" & 
    "0000011110000110" & 
    "1110000010001111" & 
    "0000000111111011" & 
    "1101110000111000" & 
    "1111110100001111" & 
    "1111011111100101" & 
    "0000011011100111" & 
    "0001100011000100" & 
    "0000110110011100" & 
    "0010000101010000" & 
    "0001011100101111" & 
    "1110101110110000" & 
    "1111101011111110" & 
    "1100111110011001" & 
    "1111011111110111" & 
    "0000101000011001" & 
    "1110101010011010" & 
    "0001001000101100" & 
    "0000100010010100" & 
    "0010001001000100" & 
    "1111110111000101" & 
    "0000000111101011" & 
    "0001100000010100" & 
    "1110110110100100" & 
    "0000100100001000" & 
    "1111000000111110" & 
    "1101010111110110" & 
    "0000011101111001" & 
    "1111001110011010" & 
    "0000001001111000" & 
    "0001101001000001" & 
    "1110100011001010" & 
    "0000111011001101" & 
    "1100111111101100" & 
    "0001010111011100" & 
    "1111011000011000" & 
    "1110100000110001" & 
    "0001001100110100" & 
    "1110010000000000" & 
    "1110111100000101" & 
    "1110110100101100" & 
    "1110110000110110" & 
    "0001111010010111" & 
    "1110011001110110" & 
    "0001001101011001" & 
    "0010000011110110" & 
    "1110011111111101" & 
    "0001111110100111" & 
    "1111101011111101" & 
    "1110110010100010" & 
    "1101110111111111" & 
    "1110101000011101" & 
    "0000111111111101" & 
    "1111010110000010" & 
    "0001001000101000" & 
    "1111101010011010" & 
    "0000101001101011" & 
    "0001011010111000" & 
    "1111100000011000" & 
    "1111010010100000" & 
    "0001011110001101" & 
    "1110111100001011" & 
    "0001001100011101" & 
    "1111101101011100" & 
    "1110001111011111" & 
    "0000010100001001" & 
    "1110111111011010" & 
    "0010001110010011" & 
    "0001000001110001" & 
    "0010000110010010" & 
    "0000011101011100" & 
    "1111110010110010" & 
    "0001100100101100" & 
    "0010001010011000" & 
    "0000111001011111" & 
    "0001101100110011" & 
    "1110100111010000" & 
    "0000011001110010" & 
    "1111011000001110" & 
    "1111110110000001" & 
    "0010000101100010" & 
    "1111111010001110" & 
    "0000101000000110" & 
    "0000111100000011" & 
    "1111010001101100" & 
    "1110100001110001" & 
    "1111000011011100" & 
    "1111001111010111" & 
    "1101010010011100" & 
    "1111001101111010" & 
    "1111001011101100" & 
    "1110110001111110" & 
    "0001100101001100" & 
    "1110110000000110" & 
    "0000000011011011" & 
    "1111001011011010" & 
    "1111100001111010" & 
    "0001111110010011" & 
    "1110010011010010" & 
    "0000001011000100" & 
    "1111111010110110" & 
    "1111001100001001" & 
    "0001001011100011" & 
    "1110000100111001" & 
    "1111100000111101" & 
    "0000111001001011" & 
    "1111011001110000" & 
    "0011011100111110" & 
    "0001011100100111" & 
    "0000111100001010" & 
    "1111111100011101" & 
    "1111010001101011" & 
    "1111100010001110" & 
    "1110000100101110" & 
    "1110110110010101" & 
    "1111110001101111" & 
    "0000001000011100" & 
    "0010000011010011" & 
    "0001000100000100" & 
    "0000010111001110" & 
    "0001011101010010" & 
    "1110111011111100" & 
    "0001101100011010" & 
    "1111010101000101" & 
    "0000111101111101" & 
    "0000011110101000" & 
    "1110110110100010" & 
    "1111101011111001" & 
    "1110010010100001" & 
    "1110010100100000" & 
    "0000011001011000" & 
    "1110100001000010" & 
    "0010111011100001" & 
    "0000111110000010" & 
    "0000111110111011" & 
    "1111111111100101" & 
    "1110111010001000" & 
    "0001110010111101" & 
    "1111100011000101" & 
    "1110111011100101" & 
    "1111110101110001" & 
    "1101111000100001" & 
    "0001101101011011" & 
    "0000101010001011" & 
    "0010001011011000" & 
    "1111101111110001" & 
    "0000011011001011" & 
    "0000011100011110" & 
    "1110101000001000" & 
    "0000011101011011" & 
    "1111101011010111" & 
    "1110000010010000" & 
    "0000110011000011" & 
    "0000011001100101" & 
    "1111101111111001" & 
    "1111011111101010" & 
    "1110111001111011" & 
    "0001000011100100" & 
    "1111011001010110" & 
    "0001011010111111" & 
    "1110010010010100" & 
    "1111000000000101" & 
    "1111011010011010" & 
    "1111010011000110" & 
    "1110100001100001" & 
    "1111101011011110" & 
    "1110000100001110" & 
    "0000101000001010" & 
    "1111101010001111" & 
    "0001000011001000" & 
    "0000110000001011" & 
    "0001000011000110" & 
    "0001110110111111" & 
    "0000110110111101" & 
    "1111011001001111" & 
    "0000011100100010" & 
    "1100000110011000" & 
    "0000110101000101" & 
    "1111001000110000" & 
    "1111111111110110" & 
    "0001100010100101" & 
    "0000111100011110" & 
    "0011000010001010" & 
    "0000011111001011" & 
    "0001011100100010" & 
    "1111101100101010" & 
    "1101101010111000" & 
    "1111111011000110" & 
    "1110011000101011" & 
    "0000010101001000" & 
    "1110111000011001" & 
    "1110100000111010" & 
    "0100010010001001" & 
    "1111010011000010" & 
    "0011001100101011" & 
    "0010001111010010" & 
    "1111010111001011" & 
    "0001001100111101" & 
    "1110110010011101" & 
    "0000001001010010" & 
    "0000101111101011" & 
    "1100100011111010" & 
    "0010001101101111" & 
    "1111100010110000" & 
    "1111110100101011" & 
    "0000101110000000" & 
    "0000010111011111" & 
    "0010010010111101" & 
    "0001010001001010" & 
    "0001111011110110" & 
    "0000000000110110" & 
    "1110101000101010" & 
    "0000111011001100" & 
    "1110010100011011" & 
    "0000100001000000" & 
    "1110111111000010" & 
    "1111011110011011" & 
    "0001100110001111" & 
    "0001010011111101" & 
    "1111111011101010" & 
    "0001010001110100" & 
    "1111111110010011" & 
    "1110111101111001" & 
    "0000010000000111" & 
    "0010011110110001" & 
    "1111001001011010" & 
    "1110011111000110" & 
    "1111101110011111" & 
    "1111001001100100" & 
    "1111111111011111" & 
    "0000101111100100" & 
    "0001101011111000" & 
    "0001001001110010" & 
    "1111011111011101" & 
    "0000110001001110" & 
    "0000001111010100" & 
    "0000001101000110" & 
    "0010001110001110" & 
    "1101001110001000" & 
    "1110101111010000" & 
    "0000001100010011" & 
    "1110100111110111" & 
    "0011010011010100" & 
    "0001100011100101" & 
    "0001110101100011" & 
    "0001110101110110" & 
    "1111100101001110" & 
    "0010000100101010" & 
    "0000001000011001" & 
    "1111110100000011" & 
    "0001010011101011" & 
    "1110110111101001" & 
    "0000000101001011" & 
    "1111001000101110" & 
    "0001011101111111" & 
    "0000011100100110" & 
    "1111111110110110" & 
    "0100010111111001" & 
    "1111100101111110" & 
    "0001110010101001" & 
    "0001001100001010" & 
    "0000010110101011" & 
    "0000101101111001" & 
    "1011101110111101" & 
    "1110100001101101" & 
    "0000001011101111" & 
    "1111010000101111" & 
    "0011010001011000" & 
    "0001010100111000" & 
    "0001110001100100" & 
    "0001010111000100" & 
    "1110010111110010" & 
    "0011001011000001" & 
    "1111001000110100" & 
    "1110001000000010" & 
    "1111110100000000" & 
    "1110010011010100" & 
    "1111100111101110" & 
    "1111010000100010" & 
    "1111101010100001" & 
    "1111011111110011" & 
    "1110010100000010" & 
    "0001101000101110" & 
    "1111011100001011" & 
    "0001010010001111" & 
    "1110110111101000" & 
    "1110100011101001" & 
    "1110101011111001" & 
    "0000000000100011" & 
    "1111010000110010" & 
    "0000111001011101" & 
    "1111011111111010" & 
    "0010001101111011" & 
    "1110110001000000" & 
    "0010100010010000" & 
    "0010101110101111" & 
    "1101110101111110" & 
    "0001001000011111" & 
    "1110010110100000" & 
    "1111110101000000" & 
    "1110100001110111" & 
    "1110011110100110" & 
    "0000110010011100" & 
    "1111000000101001" & 
    "0000010000001110" & 
    "1111100011100011" & 
    "0000000111111111" & 
    "0001011110101010" & 
    "1110110010011101" & 
    "0000110010011110" & 
    "0000001010011000" & 
    "1110111101010001" & 
    "0001001011101111" & 
    "1110110001100111" & 
    "0000101011110110" & 
    "1110111100010100" & 
    "1110001000111001" & 
    "0001001101101101" & 
    "0001010011011010" & 
    "0010100101001101" & 
    "0001001001101110" & 
    "1111010100101011" & 
    "1111110010011101" & 
    "1111101011001111" & 
    "1111101100011100" & 
    "1110001100111001" & 
    "1101110111010100" & 
    "1110010111001001" & 
    "1111001100100000" & 
    "0000001100101010" & 
    "0010011110011110" & 
    "1110101101010011" & 
    "0010111110000111" & 
    "0000001101100000" & 
    "0000111011010111" & 
    "0001000101101010" & 
    "1111111101010111" & 
    "1111000111101011" & 
    "1111100001001001" & 
    "1110001010110101" & 
    "1110100110001111" & 
    "1110010101001100" & 
    "0010000010111010" & 
    "1110110110011010" & 
    "0001100111001100" & 
    "0001101100001000" & 
    "0000000100101111" & 
    "0001110111010001" & 
    "1101110101001011" & 
    "0000101011011110" & 
    "1111011111100010" & 
    "1110111011011101" & 
    "1111001101010010" & 
    "1110110100010011" & 
    "0001001111111110" & 
    "0001110110111110" & 
    "1111111110111010" & 
    "0000001001011000" & 
    "1110111110000111" & 
    "0001000100000100" & 
    "0001001010101000" & 
    "1111001110100111" & 
    "1111100101000001" & 
    "0000011100011000" & 
    "1111011100111010" & 
    "0000100010011000" & 
    "1110100101101000" & 
    "0000001100011011" & 
    "0000100110101111" & 
    "0010010100001011" & 
    "0011000110011001" & 
    "1111011001000001" & 
    "1111101011100110" & 
    "0000100111101111" & 
    "1111111011111001" & 
    "1110010000001001" & 
    "1101101000111100" & 
    "1111011000011101" & 
    "1111111011010010" & 
    "0000111101101100" & 
    "0001000101100111" & 
    "0000010011101101" & 
    "0001001011011011" & 
    "0001000011110111" & 
    "0001001100001111" & 
    "0000000111000101" & 
    "1110100101001010" & 
    "0000000101101110" & 
    "1101010011111101" & 
    "0000000111101110" & 
    "0001000100000101" & 
    "0001011110100100" & 
    "0001110100000010" & 
    "1111000110001111" & 
    "0001011110101000" & 
    "0000010001010100" & 
    "1111010011101001" & 
    "0000101001100111" & 
    "1110001010111010" & 
    "0000000011001100" & 
    "1110010000111001" & 
    "1110110111011100" & 
    "0000111111001000" & 
    "1111110011011000" & 
    "0000010110011111" & 
    "0001011101101100" & 
    "0001110111101101" & 
    "0010000011011001" & 
    "1111111000111011" & 
    "0010100111100001" & 
    "1101110111001111" & 
    "1110010011110000" & 
    "0010100111110001" & 
    "1101101110100011" & 
    "1110110100011010" & 
    "1110011100011111" & 
    "1111110010111111" & 
    "1111001100101111" & 
    "1111000111101110" & 
    "0001110110000011" & 
    "0001010001101011" & 
    "0000100010110100" & 
    "0001011011111000" & 
    "1111101011110100" & 
    "1110011000100110" & 
    "1111100110001111" & 
    "1100101000011110" & 
    "0000111110010111" & 
    "1110011101000110" & 
    "0001000001101111" & 
    "0000010011101011" & 
    "0000011001010110" & 
    "0011000011011101" & 
    "1110000101100111" & 
    "1110111110100100" & 
    "1110100010100010" & 
    "1111100111010010" & 
    "0000100110001010" & 
    "1101011111110001" & 
    "0000111000001101" & 
    "1111110011110011" & 
    "1101011010101011" & 
    "0000010010100011" & 
    "1110100010001110" & 
    "0010001110111000" & 
    "0000101011010011" & 
    "1110101111111000" & 
    "0000101110110110" & 
    "1110001010101101" & 
    "0000100001100101" & 
    "1111110110110101" & 
    "1110100000000101" & 
    "0000100110110101" & 
    "1110110011101110" & 
    "1111011011000100" & 
    "0001011000101111" & 
    "1111001111110000" & 
    "0000111011011001" & 
    "1110111111100100" & 
    "0001101101101110" & 
    "0001010110100101" & 
    "1101000000011010" & 
    "0000000010110000" & 
    "1110011100110111" & 
    "1110110001001101" & 
    "0000011011101100" & 
    "1111010000100001" & 
    "0001001010000000" & 
    "1111010111001101" & 
    "0001111101000110" & 
    "0010001000001000" & 
    "0000011000111010" & 
    "0001000100011100" & 
    "1111111011001011" & 
    "1110110000111100" & 
    "1111100001100001" & 
    "1111100110000110" & 
    "0000000000000101" & 
    "1101111010111110" & 
    "0010010100001011" & 
    "0000100110010001" & 
    "0000100000100100" & 
    "0001001100100100" & 
    "0000010110101110" & 
    "0001010011111101" & 
    "0000011000000110" & 
    "1111000101110110" & 
    "0001011001010100" & 
    "1100110010110111" & 
    "1111100101011011" & 
    "1101101011100011" & 
    "1111000010000011" & 
    "0011001111010101" & 
    "0000110111000111" & 
    "0001010001010101" & 
    "0000111100001000" & 
    "0000011100101100" & 
    "0010010111011011" & 
    "1111000001001011" & 
    "0001010010010101" & 
    "1110100100000100" & 
    "1100001100111000" & 
    "1111011100010110" & 
    "1110100100001110" & 
    "1111111111111100" & 
    "1111111111110110" & 
    "0001011001111001" & 
    "0000011000100100" & 
    "1111100100110101" & 
    "1111111000000010" & 
    "1111111001011101" & 
    "1110000110010110" & 
    "0000101010110110" & 
    "1101001010000110" & 
    "1110100011110000" & 
    "1111110001011101" & 
    "0000000101100111" & 
    "1111011101000110" & 
    "0001101110000100" & 
    "0000011001100011" & 
    "0001111011001110" & 
    "0000111110000011" & 
    "0010101000011101" & 
    "1110011111001000" & 
    "1111101100100010" & 
    "1111001101111000" & 
    "1101100101111110" & 
    "0000011101100111" & 
    "1111000111111011" & 
    "0000000001010000" & 
    "0000111110100011" & 
    "0010101111011011" & 
    "0001111111100001" & 
    "0000110001110001" & 
    "0000011000011110" & 
    "1111110110000001" & 
    "1110011010110110" & 
    "0000110000010111" & 
    "1101011001011011" & 
    "1101100001101100" & 
    "1111101110011001" & 
    "1110100100010011" & 
    "0001100101101101" & 
    "0000000000010011" & 
    "0010000000011100" & 
    "0010001011011011" & 
    "1110100110000010" & 
    "1111110010001101" & 
    "1111100000011001" & 
    "1111111110100110" & 
    "1110011100001011" & 
    "1111011011111011" & 
    "0000001110010101" & 
    "1110111000111000" & 
    "0000101001010101" & 
    "0001100110010110" & 
    "0001100101111000" & 
    "0001101111001111" & 
    "1110010101100011" & 
    "0001110110111100" & 
    "1111011100011011" & 
    "0000000000100100" & 
    "1111100110100000" & 
    "1111101100001100" & 
    "1110100100101100" & 
    "1110100011110010" & 
    "1111111101011110" & 
    "1111111100100011" & 
    "0000100110011100" & 
    "0001101101110010" & 
    "0001001000100110" & 
    "1111100101000001" & 
    "0011010111011111" & 
    "1110101000010001" & 
    "1111011110110100" & 
    "1110011100001100" & 
    "1101011000101011" & 
    "1111100110111000" & 
    "0000011110011000" & 
    "1111111110110100" & 
    "0000001001111010" & 
    "1111100111101000" & 
    "0010101101101110" & 
    "1110110000000110" & 
    "0001011110001101" & 
    "1111000010100110" & 
    "1110101000100110" & 
    "1110010111010011" & 
    "1110101111000010" & 
    "0000000100100111" & 
    "1110111110111111" & 
    "1111010100100100" & 
    "0001011110001101" & 
    "0001000101000100" & 
    "0001011001111111" & 
    "0010010100010011" & 
    "1111110011011010" & 
    "0000101010010010" & 
    "1110111101110011" & 
    "1111011110001110" & 
    "0000010000101101" & 
    "1110001001001001" & 
    "1111010110011001" & 
    "1110100111000100" & 
    "0001100011110111" & 
    "0000011011100001" & 
    "1111011010001010" & 
    "0010111110111110" & 
    "0000001010110010" & 
    "0000011110110111" & 
    "1111101000100001" & 
    "1101010010010001" & 
    "0000010110000010" & 
    "1101111000011100" & 
    "1111101100101100" & 
    "1110001101110001" & 
    "0000010100110101" & 
    "0001110010111101" & 
    "1110010110100111" & 
    "0010010101011011" & 
    "0000101100001010" & 
    "0000001110001110" & 
    "0001100001110101" & 
    "1110001000000010" & 
    "1100110011110111" & 
    "1111111010100011" & 
    "1101110110110110" & 
    "1111100101111101" & 
    "1111001011110010" & 
    "1111101011101010" & 
    "0001100001000010" & 
    "0000001101111110" & 
    "0001000000100100" & 
    "0000111001110111" & 
    "0001010100011100" & 
    "0001100111111100" & 
    "1101110111110110" & 
    "1111010010111011" & 
    "1110100000110010" & 
    "0000000010111110" & 
    "0000011111111111" & 
    "1111000000101001" & 
    "0001000100101100" & 
    "0000100100101010" & 
    "0011001111100000" & 
    "0010001010011000" & 
    "0000000000010010" & 
    "0000101111000001" & 
    "1111100000001110" & 
    "1111001100000000" & 
    "1111100111100010" & 
    "1110111110100010" & 
    "0001000111011000" & 
    "1111010110100111" & 
    "0001101111111111" & 
    "0010101100100011" & 
    "1110001010110111" & 
    "0000001110001011" & 
    "1111001001010000" & 
    "1110110110001101" & 
    "0000000000111100" & 
    "1110011011011100" & 
    "0000011100010000" & 
    "1110011111000011" & 
    "1110101100010111" & 
    "1110110110111100" & 
    "1111110011000001" & 
    "0000111011010101" & 
    "1110100011001000" & 
    "0001010010011011" & 
    "0001011110110101" & 
    "1111100000100101" & 
    "0001111110010000" & 
    "1111001110101100" & 
    "1111011101010111" & 
    "1111010101011101" & 
    "1110101010000011" & 
    "1111101111111110" & 
    "1101101101011101" & 
    "0000001101110110" & 
    "0000111110010101" & 
    "0000100100111010" & 
    "0001111110000101" & 
    "1111100111000010" & 
    "0001011100001111" & 
    "0000010000100010" & 
    "1111100100101000" & 
    "0000000110011110" & 
    "1110001100010101" & 
    "1111010010011001" & 
    "1110110000000001" & 
    "1110000100111010" & 
    "0000010110010001" & 
    "0001101101000111" & 
    "0001000100111101" & 
    "0010001101111101" & 
    "0000010001001110" & 
    "0011001010110001" & 
    "1111111011100100" & 
    "1110011100011101" & 
    "1111000011010101" & 
    "1111000101110011" & 
    "0000011110101011" & 
    "0001000001111101" & 
    "0000010100101111" & 
    "1111010010110000" & 
    "0000100000101111" & 
    "0001000101101001"
  );

end pkg_InputSamplesFi;
